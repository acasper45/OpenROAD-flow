# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hd__dlygate4sd2_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_hd__dlygate4sd2_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  3.220000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.055000 0.625000 1.615000 ;
    END
  END A
  PIN X
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.570000 0.255000 3.135000 0.825000 ;
        RECT 2.570000 1.495000 3.135000 2.465000 ;
        RECT 2.675000 0.825000 3.135000 1.495000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 3.220000 0.085000 ;
        RECT 0.655000  0.085000 0.925000 0.545000 ;
        RECT 2.075000  0.085000 2.400000 0.545000 ;
      LAYER mcon ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
        RECT 0.605000 -0.085000 0.775000 0.085000 ;
        RECT 1.065000 -0.085000 1.235000 0.085000 ;
        RECT 1.525000 -0.085000 1.695000 0.085000 ;
        RECT 1.985000 -0.085000 2.155000 0.085000 ;
        RECT 2.445000 -0.085000 2.615000 0.085000 ;
        RECT 2.905000 -0.085000 3.075000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.240000 3.220000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 3.220000 2.805000 ;
        RECT 0.655000 2.175000 0.925000 2.635000 ;
        RECT 2.075000 2.175000 2.400000 2.635000 ;
      LAYER mcon ;
        RECT 0.145000 2.635000 0.315000 2.805000 ;
        RECT 0.605000 2.635000 0.775000 2.805000 ;
        RECT 1.065000 2.635000 1.235000 2.805000 ;
        RECT 1.525000 2.635000 1.695000 2.805000 ;
        RECT 1.985000 2.635000 2.155000 2.805000 ;
        RECT 2.445000 2.635000 2.615000 2.805000 ;
        RECT 2.905000 2.635000 3.075000 2.805000 ;
      LAYER met1 ;
        RECT 0.000000 2.480000 3.220000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085000 0.255000 0.485000 0.715000 ;
      RECT 0.085000 0.715000 1.030000 0.885000 ;
      RECT 0.085000 1.785000 1.030000 2.005000 ;
      RECT 0.085000 2.005000 0.485000 2.465000 ;
      RECT 0.795000 0.885000 1.030000 0.995000 ;
      RECT 0.795000 0.995000 1.085000 1.325000 ;
      RECT 0.795000 1.325000 1.030000 1.785000 ;
      RECT 1.155000 0.255000 1.425000 0.585000 ;
      RECT 1.155000 2.135000 1.425000 2.465000 ;
      RECT 1.255000 0.585000 1.425000 1.055000 ;
      RECT 1.255000 1.055000 2.030000 1.615000 ;
      RECT 1.255000 1.615000 1.425000 2.135000 ;
      RECT 1.615000 0.255000 1.875000 0.715000 ;
      RECT 1.615000 0.715000 2.400000 0.885000 ;
      RECT 1.615000 1.785000 2.400000 2.005000 ;
      RECT 1.615000 2.005000 1.875000 2.465000 ;
      RECT 2.200000 0.885000 2.400000 0.995000 ;
      RECT 2.200000 0.995000 2.505000 1.325000 ;
      RECT 2.200000 1.325000 2.400000 1.785000 ;
  END
END sky130_fd_sc_hd__dlygate4sd2_1
END LIBRARY
