# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hd__mux2i_4
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_hd__mux2i_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  8.280000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A0
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.560000 0.995000 1.070000 1.105000 ;
        RECT 0.560000 1.105000 1.240000 1.325000 ;
    END
  END A0
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.955000 0.995000 3.550000 1.325000 ;
    END
  END A1
  PIN S
    ANTENNAGATEAREA  1.237500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.845000 1.075000 5.930000 1.290000 ;
        RECT 5.760000 1.290000 5.930000 1.425000 ;
        RECT 5.760000 1.425000 7.850000 1.595000 ;
        RECT 7.680000 0.995000 7.850000 1.425000 ;
    END
  END S
  PIN Y
    ANTENNADIFFAREA  2.194500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.095000 0.315000 3.785000 0.485000 ;
        RECT 0.095000 0.485000 0.320000 2.255000 ;
        RECT 0.095000 2.255000 3.785000 2.425000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 8.280000 0.085000 ;
        RECT 3.975000  0.085000 4.305000 0.465000 ;
        RECT 4.815000  0.085000 5.145000 0.465000 ;
        RECT 5.655000  0.085000 5.980000 0.590000 ;
        RECT 6.545000  0.085000 6.795000 0.545000 ;
        RECT 7.435000  0.085000 7.765000 0.465000 ;
      LAYER mcon ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
        RECT 0.605000 -0.085000 0.775000 0.085000 ;
        RECT 1.065000 -0.085000 1.235000 0.085000 ;
        RECT 1.525000 -0.085000 1.695000 0.085000 ;
        RECT 1.985000 -0.085000 2.155000 0.085000 ;
        RECT 2.445000 -0.085000 2.615000 0.085000 ;
        RECT 2.905000 -0.085000 3.075000 0.085000 ;
        RECT 3.365000 -0.085000 3.535000 0.085000 ;
        RECT 3.825000 -0.085000 3.995000 0.085000 ;
        RECT 4.285000 -0.085000 4.455000 0.085000 ;
        RECT 4.745000 -0.085000 4.915000 0.085000 ;
        RECT 5.205000 -0.085000 5.375000 0.085000 ;
        RECT 5.665000 -0.085000 5.835000 0.085000 ;
        RECT 6.125000 -0.085000 6.295000 0.085000 ;
        RECT 6.585000 -0.085000 6.755000 0.085000 ;
        RECT 7.045000 -0.085000 7.215000 0.085000 ;
        RECT 7.505000 -0.085000 7.675000 0.085000 ;
        RECT 7.965000 -0.085000 8.135000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.240000 8.280000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 8.280000 2.805000 ;
        RECT 3.975000 2.255000 4.305000 2.635000 ;
        RECT 4.815000 2.255000 5.145000 2.635000 ;
        RECT 5.655000 2.255000 5.985000 2.635000 ;
        RECT 6.495000 2.255000 6.825000 2.635000 ;
        RECT 7.435000 2.255000 7.765000 2.635000 ;
      LAYER mcon ;
        RECT 0.145000 2.635000 0.315000 2.805000 ;
        RECT 0.605000 2.635000 0.775000 2.805000 ;
        RECT 1.065000 2.635000 1.235000 2.805000 ;
        RECT 1.525000 2.635000 1.695000 2.805000 ;
        RECT 1.985000 2.635000 2.155000 2.805000 ;
        RECT 2.445000 2.635000 2.615000 2.805000 ;
        RECT 2.905000 2.635000 3.075000 2.805000 ;
        RECT 3.365000 2.635000 3.535000 2.805000 ;
        RECT 3.825000 2.635000 3.995000 2.805000 ;
        RECT 4.285000 2.635000 4.455000 2.805000 ;
        RECT 4.745000 2.635000 4.915000 2.805000 ;
        RECT 5.205000 2.635000 5.375000 2.805000 ;
        RECT 5.665000 2.635000 5.835000 2.805000 ;
        RECT 6.125000 2.635000 6.295000 2.805000 ;
        RECT 6.585000 2.635000 6.755000 2.805000 ;
        RECT 7.045000 2.635000 7.215000 2.805000 ;
        RECT 7.505000 2.635000 7.675000 2.805000 ;
        RECT 7.965000 2.635000 8.135000 2.805000 ;
      LAYER met1 ;
        RECT 0.000000 2.480000 8.280000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.515000 0.655000 1.700000 0.825000 ;
      RECT 0.515000 1.575000 5.580000 1.745000 ;
      RECT 1.355000 0.825000 1.700000 0.935000 ;
      RECT 2.195000 0.655000 5.485000 0.825000 ;
      RECT 2.195000 1.915000 7.165000 2.085000 ;
      RECT 4.475000 0.255000 4.645000 0.655000 ;
      RECT 5.315000 0.255000 5.485000 0.655000 ;
      RECT 6.150000 0.255000 6.325000 0.715000 ;
      RECT 6.150000 0.715000 7.165000 0.905000 ;
      RECT 6.150000 0.905000 6.450000 0.935000 ;
      RECT 6.155000 1.795000 6.325000 1.915000 ;
      RECT 6.155000 2.085000 6.325000 2.465000 ;
      RECT 6.730000 1.075000 7.510000 1.245000 ;
      RECT 6.995000 0.510000 7.165000 0.715000 ;
      RECT 6.995000 1.795000 7.165000 1.915000 ;
      RECT 6.995000 2.085000 7.165000 2.465000 ;
      RECT 7.340000 0.655000 8.195000 0.825000 ;
      RECT 7.340000 0.825000 7.510000 1.075000 ;
      RECT 7.935000 0.255000 8.195000 0.655000 ;
      RECT 7.935000 1.795000 8.195000 2.465000 ;
      RECT 8.020000 0.825000 8.195000 1.795000 ;
    LAYER mcon ;
      RECT 1.530000 0.765000 1.700000 0.935000 ;
      RECT 6.150000 0.765000 6.320000 0.935000 ;
    LAYER met1 ;
      RECT 1.470000 0.735000 1.760000 0.780000 ;
      RECT 1.470000 0.780000 6.380000 0.920000 ;
      RECT 1.470000 0.920000 1.760000 0.965000 ;
      RECT 6.090000 0.735000 6.380000 0.780000 ;
      RECT 6.090000 0.920000 6.380000 0.965000 ;
  END
END sky130_fd_sc_hd__mux2i_4
END LIBRARY
