# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hd__nor4bb_4
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_hd__nor4bb_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.200000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.375000 1.075000 9.110000 1.285000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.150000 1.075000 7.105000 1.285000 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.110000 1.075000 0.445000 1.365000 ;
    END
  END C_N
  PIN D_N
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.955000 1.075000 1.295000 1.325000 ;
    END
  END D_N
  PIN Y
    ANTENNADIFFAREA  1.944000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.840000 1.415000 3.185000 1.705000 ;
        RECT 1.935000 0.255000 2.265000 0.725000 ;
        RECT 1.935000 0.725000 8.665000 0.905000 ;
        RECT 2.775000 0.255000 3.105000 0.725000 ;
        RECT 3.015000 0.905000 3.185000 1.415000 ;
        RECT 3.615000 0.255000 3.945000 0.725000 ;
        RECT 4.455000 0.255000 4.785000 0.725000 ;
        RECT 5.815000 0.255000 6.145000 0.725000 ;
        RECT 6.655000 0.255000 6.985000 0.725000 ;
        RECT 7.495000 0.255000 7.825000 0.725000 ;
        RECT 8.335000 0.255000 8.665000 0.725000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 9.200000 0.085000 ;
        RECT 0.615000  0.085000 0.785000 0.555000 ;
        RECT 1.595000  0.085000 1.765000 0.555000 ;
        RECT 2.435000  0.085000 2.605000 0.555000 ;
        RECT 3.275000  0.085000 3.445000 0.555000 ;
        RECT 4.115000  0.085000 4.285000 0.555000 ;
        RECT 4.955000  0.085000 5.645000 0.555000 ;
        RECT 6.315000  0.085000 6.485000 0.555000 ;
        RECT 7.155000  0.085000 7.325000 0.555000 ;
        RECT 7.995000  0.085000 8.165000 0.555000 ;
        RECT 8.835000  0.085000 9.110000 0.905000 ;
      LAYER mcon ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
        RECT 0.605000 -0.085000 0.775000 0.085000 ;
        RECT 1.065000 -0.085000 1.235000 0.085000 ;
        RECT 1.525000 -0.085000 1.695000 0.085000 ;
        RECT 1.985000 -0.085000 2.155000 0.085000 ;
        RECT 2.445000 -0.085000 2.615000 0.085000 ;
        RECT 2.905000 -0.085000 3.075000 0.085000 ;
        RECT 3.365000 -0.085000 3.535000 0.085000 ;
        RECT 3.825000 -0.085000 3.995000 0.085000 ;
        RECT 4.285000 -0.085000 4.455000 0.085000 ;
        RECT 4.745000 -0.085000 4.915000 0.085000 ;
        RECT 5.205000 -0.085000 5.375000 0.085000 ;
        RECT 5.665000 -0.085000 5.835000 0.085000 ;
        RECT 6.125000 -0.085000 6.295000 0.085000 ;
        RECT 6.585000 -0.085000 6.755000 0.085000 ;
        RECT 7.045000 -0.085000 7.215000 0.085000 ;
        RECT 7.505000 -0.085000 7.675000 0.085000 ;
        RECT 7.965000 -0.085000 8.135000 0.085000 ;
        RECT 8.425000 -0.085000 8.595000 0.085000 ;
        RECT 8.885000 -0.085000 9.055000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.240000 9.200000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 9.200000 2.805000 ;
        RECT 0.535000 2.215000 0.865000 2.635000 ;
        RECT 7.535000 1.795000 7.785000 2.635000 ;
        RECT 8.375000 1.795000 8.625000 2.635000 ;
      LAYER mcon ;
        RECT 0.145000 2.635000 0.315000 2.805000 ;
        RECT 0.605000 2.635000 0.775000 2.805000 ;
        RECT 1.065000 2.635000 1.235000 2.805000 ;
        RECT 1.525000 2.635000 1.695000 2.805000 ;
        RECT 1.985000 2.635000 2.155000 2.805000 ;
        RECT 2.445000 2.635000 2.615000 2.805000 ;
        RECT 2.905000 2.635000 3.075000 2.805000 ;
        RECT 3.365000 2.635000 3.535000 2.805000 ;
        RECT 3.825000 2.635000 3.995000 2.805000 ;
        RECT 4.285000 2.635000 4.455000 2.805000 ;
        RECT 4.745000 2.635000 4.915000 2.805000 ;
        RECT 5.205000 2.635000 5.375000 2.805000 ;
        RECT 5.665000 2.635000 5.835000 2.805000 ;
        RECT 6.125000 2.635000 6.295000 2.805000 ;
        RECT 6.585000 2.635000 6.755000 2.805000 ;
        RECT 7.045000 2.635000 7.215000 2.805000 ;
        RECT 7.505000 2.635000 7.675000 2.805000 ;
        RECT 7.965000 2.635000 8.135000 2.805000 ;
        RECT 8.425000 2.635000 8.595000 2.805000 ;
        RECT 8.885000 2.635000 9.055000 2.805000 ;
      LAYER met1 ;
        RECT 0.000000 2.480000 9.200000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.085000 0.255000 0.445000 0.725000 ;
      RECT 0.085000 0.725000 0.785000 0.895000 ;
      RECT 0.085000 1.535000 0.785000 1.875000 ;
      RECT 0.085000 1.875000 3.525000 2.045000 ;
      RECT 0.085000 2.045000 0.365000 2.465000 ;
      RECT 0.615000 0.895000 0.785000 1.535000 ;
      RECT 0.955000 0.255000 1.285000 0.735000 ;
      RECT 0.955000 0.735000 1.635000 0.905000 ;
      RECT 0.955000 1.535000 1.635000 1.705000 ;
      RECT 1.465000 0.905000 1.635000 1.075000 ;
      RECT 1.465000 1.075000 2.845000 1.245000 ;
      RECT 1.465000 1.245000 1.635000 1.535000 ;
      RECT 1.515000 2.215000 3.525000 2.295000 ;
      RECT 1.515000 2.295000 5.195000 2.465000 ;
      RECT 3.355000 1.075000 4.905000 1.285000 ;
      RECT 3.355000 1.285000 3.525000 1.875000 ;
      RECT 3.695000 1.455000 6.945000 1.625000 ;
      RECT 3.695000 1.625000 3.905000 2.125000 ;
      RECT 4.075000 1.795000 4.325000 2.295000 ;
      RECT 4.495000 1.625000 4.745000 2.125000 ;
      RECT 4.915000 1.795000 5.195000 2.295000 ;
      RECT 5.380000 1.795000 5.685000 2.295000 ;
      RECT 5.380000 2.295000 7.365000 2.465000 ;
      RECT 5.855000 1.625000 6.105000 2.125000 ;
      RECT 6.275000 1.795000 6.525000 2.295000 ;
      RECT 6.695000 1.625000 6.945000 2.125000 ;
      RECT 7.115000 1.455000 9.110000 1.625000 ;
      RECT 7.115000 1.625000 7.365000 2.295000 ;
      RECT 7.955000 1.625000 8.205000 2.465000 ;
      RECT 8.795000 1.625000 9.110000 2.465000 ;
  END
END sky130_fd_sc_hd__nor4bb_4
END LIBRARY
