# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hd__sedfxtp_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_hd__sedfxtp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  13.34000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.695000 0.765000 1.915000 1.720000 ;
    END
  END D
  PIN DE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.110000 0.765000 2.565000 1.185000 ;
        RECT 2.110000 1.185000 2.325000 1.370000 ;
    END
  END DE
  PIN Q
    ANTENNADIFFAREA  0.462000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.765000 0.305000 13.095000 2.420000 ;
    END
  END Q
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.760000 1.105000 6.215000 1.665000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 5.025000 1.105000 5.250000 1.615000 ;
    END
  END SCE
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.095000 0.975000 0.445000 1.625000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT  0.000000 -0.085000 13.340000 0.085000 ;
        RECT  0.515000  0.085000  0.845000 0.465000 ;
        RECT  2.235000  0.085000  2.565000 0.515000 ;
        RECT  3.185000  0.085000  3.515000 0.610000 ;
        RECT  5.760000  0.085000  6.010000 0.905000 ;
        RECT  8.245000  0.085000  8.640000 0.560000 ;
        RECT  9.465000  0.085000  9.740000 0.615000 ;
        RECT 11.350000  0.085000 11.665000 0.615000 ;
        RECT 12.350000  0.085000 12.595000 0.900000 ;
      LAYER mcon ;
        RECT  0.145000 -0.085000  0.315000 0.085000 ;
        RECT  0.605000 -0.085000  0.775000 0.085000 ;
        RECT  1.065000 -0.085000  1.235000 0.085000 ;
        RECT  1.525000 -0.085000  1.695000 0.085000 ;
        RECT  1.985000 -0.085000  2.155000 0.085000 ;
        RECT  2.445000 -0.085000  2.615000 0.085000 ;
        RECT  2.905000 -0.085000  3.075000 0.085000 ;
        RECT  3.365000 -0.085000  3.535000 0.085000 ;
        RECT  3.825000 -0.085000  3.995000 0.085000 ;
        RECT  4.285000 -0.085000  4.455000 0.085000 ;
        RECT  4.745000 -0.085000  4.915000 0.085000 ;
        RECT  5.205000 -0.085000  5.375000 0.085000 ;
        RECT  5.665000 -0.085000  5.835000 0.085000 ;
        RECT  6.125000 -0.085000  6.295000 0.085000 ;
        RECT  6.585000 -0.085000  6.755000 0.085000 ;
        RECT  7.045000 -0.085000  7.215000 0.085000 ;
        RECT  7.505000 -0.085000  7.675000 0.085000 ;
        RECT  7.965000 -0.085000  8.135000 0.085000 ;
        RECT  8.425000 -0.085000  8.595000 0.085000 ;
        RECT  8.885000 -0.085000  9.055000 0.085000 ;
        RECT  9.345000 -0.085000  9.515000 0.085000 ;
        RECT  9.805000 -0.085000  9.975000 0.085000 ;
        RECT 10.265000 -0.085000 10.435000 0.085000 ;
        RECT 10.725000 -0.085000 10.895000 0.085000 ;
        RECT 11.185000 -0.085000 11.355000 0.085000 ;
        RECT 11.645000 -0.085000 11.815000 0.085000 ;
        RECT 12.105000 -0.085000 12.275000 0.085000 ;
        RECT 12.565000 -0.085000 12.735000 0.085000 ;
        RECT 13.025000 -0.085000 13.195000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.240000 13.340000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT  0.000000 2.635000 13.340000 2.805000 ;
        RECT  0.515000 2.135000  0.845000 2.635000 ;
        RECT  2.235000 1.890000  2.565000 2.635000 ;
        RECT  3.265000 1.825000  3.460000 2.635000 ;
        RECT  5.665000 2.175000  6.010000 2.635000 ;
        RECT  8.425000 1.835000  8.660000 2.635000 ;
        RECT  9.370000 2.105000  9.660000 2.635000 ;
        RECT 11.280000 2.135000 11.540000 2.635000 ;
        RECT 12.350000 1.465000 12.595000 2.635000 ;
      LAYER mcon ;
        RECT  0.145000 2.635000  0.315000 2.805000 ;
        RECT  0.605000 2.635000  0.775000 2.805000 ;
        RECT  1.065000 2.635000  1.235000 2.805000 ;
        RECT  1.525000 2.635000  1.695000 2.805000 ;
        RECT  1.985000 2.635000  2.155000 2.805000 ;
        RECT  2.445000 2.635000  2.615000 2.805000 ;
        RECT  2.905000 2.635000  3.075000 2.805000 ;
        RECT  3.365000 2.635000  3.535000 2.805000 ;
        RECT  3.825000 2.635000  3.995000 2.805000 ;
        RECT  4.285000 2.635000  4.455000 2.805000 ;
        RECT  4.745000 2.635000  4.915000 2.805000 ;
        RECT  5.205000 2.635000  5.375000 2.805000 ;
        RECT  5.665000 2.635000  5.835000 2.805000 ;
        RECT  6.125000 2.635000  6.295000 2.805000 ;
        RECT  6.585000 2.635000  6.755000 2.805000 ;
        RECT  7.045000 2.635000  7.215000 2.805000 ;
        RECT  7.505000 2.635000  7.675000 2.805000 ;
        RECT  7.965000 2.635000  8.135000 2.805000 ;
        RECT  8.425000 2.635000  8.595000 2.805000 ;
        RECT  8.885000 2.635000  9.055000 2.805000 ;
        RECT  9.345000 2.635000  9.515000 2.805000 ;
        RECT  9.805000 2.635000  9.975000 2.805000 ;
        RECT 10.265000 2.635000 10.435000 2.805000 ;
        RECT 10.725000 2.635000 10.895000 2.805000 ;
        RECT 11.185000 2.635000 11.355000 2.805000 ;
        RECT 11.645000 2.635000 11.815000 2.805000 ;
        RECT 12.105000 2.635000 12.275000 2.805000 ;
        RECT 12.565000 2.635000 12.735000 2.805000 ;
        RECT 13.025000 2.635000 13.195000 2.805000 ;
      LAYER met1 ;
        RECT 0.000000 2.480000 13.340000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.175000 0.345000  0.345000 0.635000 ;
      RECT  0.175000 0.635000  0.845000 0.805000 ;
      RECT  0.175000 1.795000  0.845000 1.965000 ;
      RECT  0.175000 1.965000  0.345000 2.465000 ;
      RECT  0.615000 0.805000  0.845000 1.795000 ;
      RECT  1.015000 0.345000  1.185000 2.465000 ;
      RECT  1.355000 0.255000  1.785000 0.515000 ;
      RECT  1.355000 0.515000  1.525000 1.890000 ;
      RECT  1.355000 1.890000  1.785000 2.465000 ;
      RECT  2.495000 1.355000  3.085000 1.720000 ;
      RECT  2.755000 1.720000  3.085000 2.425000 ;
      RECT  2.780000 0.255000  3.005000 0.845000 ;
      RECT  2.780000 0.845000  3.635000 1.175000 ;
      RECT  2.780000 1.175000  3.085000 1.355000 ;
      RECT  3.805000 0.685000  3.975000 1.320000 ;
      RECT  3.805000 1.320000  4.175000 1.650000 ;
      RECT  4.125000 1.820000  4.515000 2.020000 ;
      RECT  4.125000 2.020000  4.455000 2.465000 ;
      RECT  4.145000 0.255000  4.415000 0.980000 ;
      RECT  4.145000 0.980000  4.515000 1.150000 ;
      RECT  4.345000 1.150000  4.515000 1.820000 ;
      RECT  4.595000 0.255000  4.795000 0.645000 ;
      RECT  4.595000 0.645000  4.855000 0.825000 ;
      RECT  4.635000 2.210000  4.965000 2.465000 ;
      RECT  4.685000 0.825000  4.855000 1.785000 ;
      RECT  4.685000 1.785000  4.965000 2.210000 ;
      RECT  4.965000 0.255000  5.590000 0.515000 ;
      RECT  5.155000 1.835000  6.585000 2.005000 ;
      RECT  5.155000 2.005000  5.495000 2.465000 ;
      RECT  5.260000 0.515000  5.590000 0.935000 ;
      RECT  5.420000 0.935000  5.590000 1.835000 ;
      RECT  6.385000 1.355000  6.585000 1.835000 ;
      RECT  6.515000 0.255000  7.135000 0.565000 ;
      RECT  6.515000 0.565000  6.925000 1.185000 ;
      RECT  6.675000 2.150000  7.005000 2.465000 ;
      RECT  6.755000 1.185000  6.925000 1.865000 ;
      RECT  6.755000 1.865000  7.005000 2.150000 ;
      RECT  7.095000 1.125000  7.280000 1.720000 ;
      RECT  7.115000 0.735000  7.620000 0.955000 ;
      RECT  7.215000 2.175000  8.255000 2.375000 ;
      RECT  7.305000 0.255000  7.980000 0.565000 ;
      RECT  7.450000 0.955000  7.620000 1.655000 ;
      RECT  7.450000 1.655000  7.915000 2.005000 ;
      RECT  7.810000 0.565000  7.980000 1.315000 ;
      RECT  7.810000 1.315000  8.660000 1.485000 ;
      RECT  8.085000 1.485000  8.660000 1.575000 ;
      RECT  8.085000 1.575000  8.255000 2.175000 ;
      RECT  8.170000 0.765000  9.235000 1.045000 ;
      RECT  8.170000 1.045000  9.745000 1.065000 ;
      RECT  8.170000 1.065000  8.370000 1.095000 ;
      RECT  8.490000 1.245000  8.660000 1.315000 ;
      RECT  8.830000 0.255000  9.235000 0.765000 ;
      RECT  8.830000 1.065000  9.745000 1.375000 ;
      RECT  8.830000 1.375000  9.160000 2.465000 ;
      RECT 10.090000 1.245000 10.280000 1.965000 ;
      RECT 10.225000 2.165000 11.110000 2.355000 ;
      RECT 10.305000 0.705000 10.770000 1.035000 ;
      RECT 10.325000 0.330000 11.110000 0.535000 ;
      RECT 10.450000 1.035000 10.770000 1.995000 ;
      RECT 10.940000 0.535000 11.110000 0.995000 ;
      RECT 10.940000 0.995000 11.810000 1.325000 ;
      RECT 10.940000 1.325000 11.110000 2.165000 ;
      RECT 11.280000 1.530000 12.180000 1.905000 ;
      RECT 11.840000 1.905000 12.180000 2.465000 ;
      RECT 11.850000 0.300000 12.180000 0.825000 ;
      RECT 11.990000 0.825000 12.180000 1.530000 ;
    LAYER mcon ;
      RECT  0.635000 1.785000  0.805000 1.955000 ;
      RECT  1.015000 1.445000  1.185000 1.615000 ;
      RECT  1.355000 0.425000  1.525000 0.595000 ;
      RECT  3.805000 0.765000  3.975000 0.935000 ;
      RECT  4.185000 0.425000  4.355000 0.595000 ;
      RECT  4.615000 0.425000  4.785000 0.595000 ;
      RECT  6.530000 0.425000  6.700000 0.595000 ;
      RECT  7.100000 1.445000  7.270000 1.615000 ;
      RECT  7.510000 1.785000  7.680000 1.955000 ;
      RECT 10.100000 1.785000 10.270000 1.955000 ;
      RECT 10.520000 1.445000 10.690000 1.615000 ;
      RECT 12.000000 0.765000 12.170000 0.935000 ;
    LAYER met1 ;
      RECT  0.575000 1.755000  0.865000 1.800000 ;
      RECT  0.575000 1.800000 10.330000 1.940000 ;
      RECT  0.575000 1.940000  0.865000 1.985000 ;
      RECT  0.955000 1.415000  1.245000 1.460000 ;
      RECT  0.955000 1.460000 10.750000 1.600000 ;
      RECT  0.955000 1.600000  1.245000 1.645000 ;
      RECT  1.295000 0.395000  4.415000 0.580000 ;
      RECT  1.295000 0.580000  1.585000 0.625000 ;
      RECT  3.745000 0.735000  4.035000 0.780000 ;
      RECT  3.745000 0.780000 12.230000 0.920000 ;
      RECT  3.745000 0.920000  4.035000 0.965000 ;
      RECT  4.125000 0.580000  4.415000 0.625000 ;
      RECT  4.555000 0.395000  6.760000 0.580000 ;
      RECT  4.555000 0.580000  4.845000 0.625000 ;
      RECT  6.470000 0.580000  6.760000 0.625000 ;
      RECT  7.040000 1.415000  7.330000 1.460000 ;
      RECT  7.040000 1.600000  7.330000 1.645000 ;
      RECT  7.450000 1.755000  7.740000 1.800000 ;
      RECT  7.450000 1.940000  7.740000 1.985000 ;
      RECT 10.040000 1.755000 10.330000 1.800000 ;
      RECT 10.040000 1.940000 10.330000 1.985000 ;
      RECT 10.460000 1.415000 10.750000 1.460000 ;
      RECT 10.460000 1.600000 10.750000 1.645000 ;
      RECT 11.940000 0.735000 12.230000 0.780000 ;
      RECT 11.940000 0.920000 12.230000 0.965000 ;
  END
END sky130_fd_sc_hd__sedfxtp_1
END LIBRARY
