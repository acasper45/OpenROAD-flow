# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hd__o31ai_4
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_hd__o31ai_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  7.820000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.090000 1.055000 1.780000 1.425000 ;
    END
  END A1
  PIN A2
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.950000 1.055000 3.605000 1.425000 ;
    END
  END A2
  PIN A3
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.775000 1.055000 5.940000 1.275000 ;
    END
  END A3
  PIN B1
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.465000 1.055000 7.735000 1.275000 ;
    END
  END B1
  PIN Y
    ANTENNADIFFAREA  1.683800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.775000 1.445000 7.735000 1.695000 ;
        RECT 5.770000 1.695000 5.940000 2.465000 ;
        RECT 6.110000 0.645000 7.280000 0.885000 ;
        RECT 6.110000 0.885000 6.295000 1.445000 ;
        RECT 6.610000 1.695000 6.780000 2.465000 ;
        RECT 7.450000 1.695000 7.735000 2.465000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 7.820000 0.085000 ;
        RECT 0.615000  0.085000 0.785000 0.545000 ;
        RECT 1.455000  0.085000 1.625000 0.545000 ;
        RECT 2.295000  0.085000 2.465000 0.545000 ;
        RECT 3.135000  0.085000 3.305000 0.545000 ;
        RECT 3.995000  0.085000 4.640000 0.545000 ;
        RECT 5.150000  0.085000 5.600000 0.545000 ;
      LAYER mcon ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
        RECT 0.605000 -0.085000 0.775000 0.085000 ;
        RECT 1.065000 -0.085000 1.235000 0.085000 ;
        RECT 1.525000 -0.085000 1.695000 0.085000 ;
        RECT 1.985000 -0.085000 2.155000 0.085000 ;
        RECT 2.445000 -0.085000 2.615000 0.085000 ;
        RECT 2.905000 -0.085000 3.075000 0.085000 ;
        RECT 3.365000 -0.085000 3.535000 0.085000 ;
        RECT 3.825000 -0.085000 3.995000 0.085000 ;
        RECT 4.285000 -0.085000 4.455000 0.085000 ;
        RECT 4.745000 -0.085000 4.915000 0.085000 ;
        RECT 5.205000 -0.085000 5.375000 0.085000 ;
        RECT 5.665000 -0.085000 5.835000 0.085000 ;
        RECT 6.125000 -0.085000 6.295000 0.085000 ;
        RECT 6.585000 -0.085000 6.755000 0.085000 ;
        RECT 7.045000 -0.085000 7.215000 0.085000 ;
        RECT 7.505000 -0.085000 7.675000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.240000 7.820000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 7.820000 2.805000 ;
        RECT 0.615000 2.065000 0.785000 2.635000 ;
        RECT 1.455000 2.065000 1.625000 2.635000 ;
        RECT 6.110000 1.890000 6.440000 2.635000 ;
        RECT 6.950000 1.890000 7.280000 2.635000 ;
      LAYER mcon ;
        RECT 0.145000 2.635000 0.315000 2.805000 ;
        RECT 0.605000 2.635000 0.775000 2.805000 ;
        RECT 1.065000 2.635000 1.235000 2.805000 ;
        RECT 1.525000 2.635000 1.695000 2.805000 ;
        RECT 1.985000 2.635000 2.155000 2.805000 ;
        RECT 2.445000 2.635000 2.615000 2.805000 ;
        RECT 2.905000 2.635000 3.075000 2.805000 ;
        RECT 3.365000 2.635000 3.535000 2.805000 ;
        RECT 3.825000 2.635000 3.995000 2.805000 ;
        RECT 4.285000 2.635000 4.455000 2.805000 ;
        RECT 4.745000 2.635000 4.915000 2.805000 ;
        RECT 5.205000 2.635000 5.375000 2.805000 ;
        RECT 5.665000 2.635000 5.835000 2.805000 ;
        RECT 6.125000 2.635000 6.295000 2.805000 ;
        RECT 6.585000 2.635000 6.755000 2.805000 ;
        RECT 7.045000 2.635000 7.215000 2.805000 ;
        RECT 7.505000 2.635000 7.675000 2.805000 ;
      LAYER met1 ;
        RECT 0.000000 2.480000 7.820000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.090000 0.255000 0.445000 0.715000 ;
      RECT 0.090000 0.715000 5.940000 0.885000 ;
      RECT 0.090000 1.595000 2.125000 1.895000 ;
      RECT 0.090000 1.895000 0.445000 2.465000 ;
      RECT 0.955000 0.255000 1.285000 0.715000 ;
      RECT 0.955000 1.895000 1.285000 2.465000 ;
      RECT 1.795000 0.255000 2.125000 0.715000 ;
      RECT 1.795000 1.895000 2.125000 2.205000 ;
      RECT 1.795000 2.205000 3.885000 2.465000 ;
      RECT 2.295000 1.595000 3.605000 1.765000 ;
      RECT 2.295000 1.765000 2.465000 2.035000 ;
      RECT 2.635000 0.255000 2.965000 0.715000 ;
      RECT 2.635000 1.935000 2.965000 2.205000 ;
      RECT 3.135000 1.765000 3.605000 1.865000 ;
      RECT 3.135000 1.865000 5.600000 2.035000 ;
      RECT 3.475000 0.255000 3.805000 0.715000 ;
      RECT 4.080000 2.035000 5.600000 2.465000 ;
      RECT 4.810000 0.395000 4.980000 0.715000 ;
      RECT 5.770000 0.255000 7.735000 0.475000 ;
      RECT 5.770000 0.475000 5.940000 0.715000 ;
      RECT 7.450000 0.475000 7.735000 0.885000 ;
  END
END sky130_fd_sc_hd__o31ai_4
END LIBRARY
