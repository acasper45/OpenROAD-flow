# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hd__sdfstp_4
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_hd__sdfstp_4 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  13.80000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.050000 0.765000 1.335000 1.675000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.891000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 12.040000 0.275000 12.370000 0.825000 ;
        RECT 12.040000 1.495000 12.370000 2.450000 ;
        RECT 12.145000 0.825000 12.370000 1.055000 ;
        RECT 12.145000 1.055000 13.210000 1.325000 ;
        RECT 12.145000 1.325000 12.370000 1.495000 ;
        RECT 12.880000 0.255000 13.210000 1.055000 ;
        RECT 12.880000 1.325000 13.210000 2.465000 ;
    END
  END Q
  PIN SCD
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 0.765000 0.340000 1.675000 ;
    END
  END SCD
  PIN SCE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.540000 0.765000 0.820000 1.675000 ;
        RECT 2.370000 1.075000 2.700000 1.600000 ;
      LAYER mcon ;
        RECT 0.605000 1.105000 0.775000 1.275000 ;
        RECT 2.445000 1.105000 2.615000 1.275000 ;
      LAYER met1 ;
        RECT 0.545000 1.075000 0.835000 1.120000 ;
        RECT 0.545000 1.120000 2.675000 1.260000 ;
        RECT 0.545000 1.260000 0.835000 1.305000 ;
        RECT 2.385000 1.075000 2.675000 1.120000 ;
        RECT 2.385000 1.260000 2.675000 1.305000 ;
    END
  END SCE
  PIN SET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 6.640000 1.445000 7.065000 1.765000 ;
        RECT 8.880000 1.425000 9.135000 1.545000 ;
        RECT 8.880000 1.545000 9.945000 1.725000 ;
      LAYER mcon ;
        RECT 8.940000 1.445000 9.110000 1.615000 ;
      LAYER met1 ;
        RECT 6.580000 1.415000 6.870000 1.460000 ;
        RECT 6.580000 1.460000 9.170000 1.600000 ;
        RECT 6.580000 1.600000 6.870000 1.645000 ;
        RECT 8.880000 1.415000 9.170000 1.460000 ;
        RECT 8.880000 1.600000 9.170000 1.645000 ;
    END
  END SET_B
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 2.905000 0.725000 3.100000 1.055000 ;
        RECT 2.905000 1.055000 3.565000 1.615000 ;
        RECT 2.905000 1.615000 3.085000 1.960000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT  0.000000 -0.085000 13.800000 0.085000 ;
        RECT  0.085000  0.085000  0.700000 0.595000 ;
        RECT  1.825000  0.085000  2.090000 0.545000 ;
        RECT  2.690000  0.085000  3.100000 0.555000 ;
        RECT  3.625000  0.085000  3.955000 0.545000 ;
        RECT  5.610000  0.085000  6.095000 0.465000 ;
        RECT  6.705000  0.085000  7.715000 0.805000 ;
        RECT 10.115000  0.085000 10.365000 0.545000 ;
        RECT 11.515000  0.085000 11.870000 0.825000 ;
        RECT 12.540000  0.085000 12.710000 0.885000 ;
        RECT 13.380000  0.085000 13.715000 0.885000 ;
      LAYER mcon ;
        RECT  0.145000 -0.085000  0.315000 0.085000 ;
        RECT  0.605000 -0.085000  0.775000 0.085000 ;
        RECT  1.065000 -0.085000  1.235000 0.085000 ;
        RECT  1.525000 -0.085000  1.695000 0.085000 ;
        RECT  1.985000 -0.085000  2.155000 0.085000 ;
        RECT  2.445000 -0.085000  2.615000 0.085000 ;
        RECT  2.905000 -0.085000  3.075000 0.085000 ;
        RECT  3.365000 -0.085000  3.535000 0.085000 ;
        RECT  3.825000 -0.085000  3.995000 0.085000 ;
        RECT  4.285000 -0.085000  4.455000 0.085000 ;
        RECT  4.745000 -0.085000  4.915000 0.085000 ;
        RECT  5.205000 -0.085000  5.375000 0.085000 ;
        RECT  5.665000 -0.085000  5.835000 0.085000 ;
        RECT  6.125000 -0.085000  6.295000 0.085000 ;
        RECT  6.585000 -0.085000  6.755000 0.085000 ;
        RECT  7.045000 -0.085000  7.215000 0.085000 ;
        RECT  7.505000 -0.085000  7.675000 0.085000 ;
        RECT  7.965000 -0.085000  8.135000 0.085000 ;
        RECT  8.425000 -0.085000  8.595000 0.085000 ;
        RECT  8.885000 -0.085000  9.055000 0.085000 ;
        RECT  9.345000 -0.085000  9.515000 0.085000 ;
        RECT  9.805000 -0.085000  9.975000 0.085000 ;
        RECT 10.265000 -0.085000 10.435000 0.085000 ;
        RECT 10.725000 -0.085000 10.895000 0.085000 ;
        RECT 11.185000 -0.085000 11.355000 0.085000 ;
        RECT 11.645000 -0.085000 11.815000 0.085000 ;
        RECT 12.105000 -0.085000 12.275000 0.085000 ;
        RECT 12.565000 -0.085000 12.735000 0.085000 ;
        RECT 13.025000 -0.085000 13.195000 0.085000 ;
        RECT 13.485000 -0.085000 13.655000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.240000 13.800000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT  0.000000 2.635000 13.800000 2.805000 ;
        RECT  0.515000 2.195000  0.785000 2.635000 ;
        RECT  2.690000 2.140000  2.985000 2.635000 ;
        RECT  3.595000 2.275000  3.925000 2.635000 ;
        RECT  5.945000 2.275000  6.330000 2.635000 ;
        RECT  7.060000 2.125000  8.015000 2.635000 ;
        RECT  9.160000 2.235000  9.490000 2.635000 ;
        RECT 10.155000 2.235000 10.485000 2.635000 ;
        RECT 11.515000 1.495000 11.870000 2.635000 ;
        RECT 12.540000 1.495000 12.710000 2.635000 ;
        RECT 13.380000 1.495000 13.715000 2.635000 ;
      LAYER mcon ;
        RECT  0.145000 2.635000  0.315000 2.805000 ;
        RECT  0.605000 2.635000  0.775000 2.805000 ;
        RECT  1.065000 2.635000  1.235000 2.805000 ;
        RECT  1.525000 2.635000  1.695000 2.805000 ;
        RECT  1.985000 2.635000  2.155000 2.805000 ;
        RECT  2.445000 2.635000  2.615000 2.805000 ;
        RECT  2.905000 2.635000  3.075000 2.805000 ;
        RECT  3.365000 2.635000  3.535000 2.805000 ;
        RECT  3.825000 2.635000  3.995000 2.805000 ;
        RECT  4.285000 2.635000  4.455000 2.805000 ;
        RECT  4.745000 2.635000  4.915000 2.805000 ;
        RECT  5.205000 2.635000  5.375000 2.805000 ;
        RECT  5.665000 2.635000  5.835000 2.805000 ;
        RECT  6.125000 2.635000  6.295000 2.805000 ;
        RECT  6.585000 2.635000  6.755000 2.805000 ;
        RECT  7.045000 2.635000  7.215000 2.805000 ;
        RECT  7.505000 2.635000  7.675000 2.805000 ;
        RECT  7.965000 2.635000  8.135000 2.805000 ;
        RECT  8.425000 2.635000  8.595000 2.805000 ;
        RECT  8.885000 2.635000  9.055000 2.805000 ;
        RECT  9.345000 2.635000  9.515000 2.805000 ;
        RECT  9.805000 2.635000  9.975000 2.805000 ;
        RECT 10.265000 2.635000 10.435000 2.805000 ;
        RECT 10.725000 2.635000 10.895000 2.805000 ;
        RECT 11.185000 2.635000 11.355000 2.805000 ;
        RECT 11.645000 2.635000 11.815000 2.805000 ;
        RECT 12.105000 2.635000 12.275000 2.805000 ;
        RECT 12.565000 2.635000 12.735000 2.805000 ;
        RECT 13.025000 2.635000 13.195000 2.805000 ;
        RECT 13.485000 2.635000 13.655000 2.805000 ;
      LAYER met1 ;
        RECT 0.000000 2.480000 13.800000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT  0.085000 1.845000  1.125000 2.025000 ;
      RECT  0.085000 2.025000  0.345000 2.465000 ;
      RECT  0.870000 0.255000  1.625000 0.555000 ;
      RECT  0.870000 0.555000  1.640000 0.575000 ;
      RECT  0.870000 0.575000  1.650000 0.595000 ;
      RECT  0.955000 2.025000  1.125000 2.255000 ;
      RECT  0.955000 2.255000  2.045000 2.465000 ;
      RECT  1.295000 1.845000  1.695000 2.085000 ;
      RECT  1.380000 0.595000  1.660000 0.600000 ;
      RECT  1.395000 0.600000  1.660000 0.605000 ;
      RECT  1.405000 0.605000  1.660000 0.610000 ;
      RECT  1.420000 0.610000  1.660000 0.615000 ;
      RECT  1.430000 0.615000  1.660000 0.620000 ;
      RECT  1.440000 0.620000  1.665000 0.630000 ;
      RECT  1.445000 0.630000  1.665000 0.635000 ;
      RECT  1.460000 0.635000  1.665000 0.645000 ;
      RECT  1.475000 0.645000  1.670000 0.660000 ;
      RECT  1.475000 0.660000  1.675000 0.665000 ;
      RECT  1.495000 0.665000  1.675000 0.705000 ;
      RECT  1.505000 0.705000  1.675000 0.710000 ;
      RECT  1.505000 0.710000  1.695000 1.845000 ;
      RECT  1.865000 0.715000  2.520000 0.905000 ;
      RECT  1.865000 0.905000  2.200000 1.770000 ;
      RECT  1.865000 1.770000  2.520000 2.085000 ;
      RECT  2.260000 0.255000  2.520000 0.715000 ;
      RECT  2.270000 2.085000  2.520000 2.465000 ;
      RECT  3.255000 1.830000  3.995000 1.990000 ;
      RECT  3.255000 1.990000  3.985000 2.000000 ;
      RECT  3.255000 2.000000  3.425000 2.325000 ;
      RECT  3.270000 0.255000  3.455000 0.715000 ;
      RECT  3.270000 0.715000  3.995000 0.885000 ;
      RECT  3.735000 0.885000  3.995000 1.830000 ;
      RECT  4.095000 2.135000  4.440000 2.465000 ;
      RECT  4.125000 0.255000  4.335000 0.585000 ;
      RECT  4.165000 0.585000  4.335000 1.090000 ;
      RECT  4.165000 1.090000  4.490000 1.420000 ;
      RECT  4.165000 1.420000  4.440000 2.135000 ;
      RECT  4.505000 0.255000  4.830000 0.920000 ;
      RECT  4.615000 1.590000  4.915000 1.615000 ;
      RECT  4.615000 1.615000  4.830000 2.465000 ;
      RECT  4.660000 0.920000  4.830000 1.445000 ;
      RECT  4.660000 1.445000  4.915000 1.590000 ;
      RECT  5.000000 0.255000  5.440000 1.225000 ;
      RECT  5.000000 1.225000  7.715000 1.275000 ;
      RECT  5.035000 2.135000  5.755000 2.465000 ;
      RECT  5.085000 1.275000  6.475000 1.395000 ;
      RECT  5.205000 1.575000  5.415000 1.955000 ;
      RECT  5.585000 1.395000  5.755000 2.135000 ;
      RECT  5.645000 0.635000  6.535000 0.805000 ;
      RECT  5.645000 0.805000  5.975000 1.015000 ;
      RECT  5.925000 1.575000  6.095000 1.935000 ;
      RECT  5.925000 1.935000  6.820000 2.105000 ;
      RECT  6.285000 0.255000  6.535000 0.635000 ;
      RECT  6.305000 0.975000  7.715000 1.225000 ;
      RECT  6.605000 2.105000  6.820000 2.450000 ;
      RECT  7.235000 1.670000  8.135000 1.955000 ;
      RECT  7.355000 1.275000  7.715000 1.325000 ;
      RECT  7.885000 0.720000  9.105000 0.905000 ;
      RECT  7.885000 0.905000  8.135000 1.670000 ;
      RECT  8.185000 2.125000  8.990000 2.460000 ;
      RECT  8.425000 1.075000  8.650000 1.905000 ;
      RECT  8.465000 0.275000  9.910000 0.545000 ;
      RECT  8.820000 0.905000  9.105000 1.255000 ;
      RECT  8.820000 1.895000 10.485000 2.065000 ;
      RECT  8.820000 2.065000  8.990000 2.125000 ;
      RECT  9.320000 0.855000  9.530000 1.195000 ;
      RECT  9.320000 1.195000 10.915000 1.365000 ;
      RECT  9.660000 2.065000  9.965000 2.450000 ;
      RECT  9.710000 0.545000  9.910000 0.785000 ;
      RECT  9.710000 0.785000 10.515000 1.015000 ;
      RECT 10.155000 1.605000 10.485000 1.895000 ;
      RECT 10.575000 0.255000 10.915000 0.585000 ;
      RECT 10.655000 1.365000 10.915000 2.465000 ;
      RECT 10.685000 0.585000 10.915000 1.195000 ;
      RECT 11.085000 0.255000 11.345000 0.995000 ;
      RECT 11.085000 0.995000 11.975000 1.325000 ;
      RECT 11.085000 1.325000 11.345000 2.465000 ;
    LAYER mcon ;
      RECT 1.525000 1.445000 1.695000 1.615000 ;
      RECT 3.825000 1.785000 3.995000 1.955000 ;
      RECT 4.285000 1.105000 4.455000 1.275000 ;
      RECT 4.745000 1.445000 4.915000 1.615000 ;
      RECT 5.205000 1.785000 5.375000 1.955000 ;
      RECT 7.560000 1.785000 7.730000 1.955000 ;
      RECT 8.480000 1.105000 8.650000 1.275000 ;
    LAYER met1 ;
      RECT 1.465000 1.415000 1.755000 1.460000 ;
      RECT 1.465000 1.460000 4.975000 1.600000 ;
      RECT 1.465000 1.600000 1.755000 1.645000 ;
      RECT 3.765000 1.755000 4.055000 1.800000 ;
      RECT 3.765000 1.800000 7.790000 1.940000 ;
      RECT 3.765000 1.940000 4.055000 1.985000 ;
      RECT 4.225000 1.075000 4.515000 1.120000 ;
      RECT 4.225000 1.120000 8.710000 1.260000 ;
      RECT 4.225000 1.260000 4.515000 1.305000 ;
      RECT 4.685000 1.415000 4.975000 1.460000 ;
      RECT 4.685000 1.600000 4.975000 1.645000 ;
      RECT 5.145000 1.755000 5.435000 1.800000 ;
      RECT 5.145000 1.940000 5.435000 1.985000 ;
      RECT 7.500000 1.755000 7.790000 1.800000 ;
      RECT 7.500000 1.940000 7.790000 1.985000 ;
      RECT 8.420000 1.075000 8.710000 1.120000 ;
      RECT 8.420000 1.260000 8.710000 1.305000 ;
  END
END sky130_fd_sc_hd__sdfstp_4
END LIBRARY
