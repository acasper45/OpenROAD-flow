# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hd__dfrbp_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_hd__dfrbp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  10.58000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.355000 1.665000 1.680000 2.450000 ;
        RECT 1.415000 0.615000 1.875000 1.665000 ;
    END
  END D
  PIN Q
    ANTENNADIFFAREA  0.449000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 8.600000 1.455000 9.005000 2.465000 ;
        RECT 8.675000 0.275000 9.005000 1.455000 ;
    END
  END Q
  PIN Q_N
    ANTENNADIFFAREA  0.429000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.180000 0.265000 10.435000 0.795000 ;
        RECT 10.180000 1.445000 10.435000 2.325000 ;
        RECT 10.225000 0.795000 10.435000 1.445000 ;
    END
  END Q_N
  PIN RESET_B
    ANTENNAGATEAREA  0.252000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.805000 0.765000 4.595000 1.015000 ;
        RECT 7.105000 1.035000 7.645000 1.405000 ;
        RECT 7.405000 0.635000 7.645000 1.035000 ;
      LAYER mcon ;
        RECT 4.165000 0.765000 4.335000 0.935000 ;
        RECT 7.105000 1.080000 7.275000 1.250000 ;
        RECT 7.405000 0.765000 7.575000 0.935000 ;
      LAYER met1 ;
        RECT 3.745000 0.735000 4.395000 0.780000 ;
        RECT 3.745000 0.780000 7.635000 0.920000 ;
        RECT 3.745000 0.920000 4.395000 0.965000 ;
        RECT 7.045000 0.920000 7.635000 0.965000 ;
        RECT 7.045000 0.965000 7.335000 1.280000 ;
        RECT 7.345000 0.735000 7.635000 0.780000 ;
    END
  END RESET_B
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.090000 0.975000 0.440000 1.625000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 10.580000 0.085000 ;
        RECT 0.515000  0.085000  0.845000 0.465000 ;
        RECT 1.545000  0.085000  1.875000 0.445000 ;
        RECT 4.475000  0.085000  4.805000 0.545000 ;
        RECT 6.705000  0.085000  6.895000 0.525000 ;
        RECT 8.335000  0.085000  8.505000 0.770000 ;
        RECT 9.760000  0.085000  9.930000 0.680000 ;
      LAYER mcon ;
        RECT  0.145000 -0.085000  0.315000 0.085000 ;
        RECT  0.605000 -0.085000  0.775000 0.085000 ;
        RECT  1.065000 -0.085000  1.235000 0.085000 ;
        RECT  1.525000 -0.085000  1.695000 0.085000 ;
        RECT  1.985000 -0.085000  2.155000 0.085000 ;
        RECT  2.445000 -0.085000  2.615000 0.085000 ;
        RECT  2.905000 -0.085000  3.075000 0.085000 ;
        RECT  3.365000 -0.085000  3.535000 0.085000 ;
        RECT  3.825000 -0.085000  3.995000 0.085000 ;
        RECT  4.285000 -0.085000  4.455000 0.085000 ;
        RECT  4.745000 -0.085000  4.915000 0.085000 ;
        RECT  5.205000 -0.085000  5.375000 0.085000 ;
        RECT  5.665000 -0.085000  5.835000 0.085000 ;
        RECT  6.125000 -0.085000  6.295000 0.085000 ;
        RECT  6.585000 -0.085000  6.755000 0.085000 ;
        RECT  7.045000 -0.085000  7.215000 0.085000 ;
        RECT  7.505000 -0.085000  7.675000 0.085000 ;
        RECT  7.965000 -0.085000  8.135000 0.085000 ;
        RECT  8.425000 -0.085000  8.595000 0.085000 ;
        RECT  8.885000 -0.085000  9.055000 0.085000 ;
        RECT  9.345000 -0.085000  9.515000 0.085000 ;
        RECT  9.805000 -0.085000  9.975000 0.085000 ;
        RECT 10.265000 -0.085000 10.435000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.240000 10.580000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 10.580000 2.805000 ;
        RECT 0.515000 2.135000  0.845000 2.635000 ;
        RECT 1.850000 2.175000  2.100000 2.635000 ;
        RECT 3.990000 2.205000  4.320000 2.635000 ;
        RECT 4.955000 2.175000  5.325000 2.635000 ;
        RECT 6.940000 2.175000  7.190000 2.635000 ;
        RECT 7.710000 2.255000  8.430000 2.635000 ;
        RECT 9.760000 1.495000  9.930000 2.635000 ;
      LAYER mcon ;
        RECT  0.145000 2.635000  0.315000 2.805000 ;
        RECT  0.605000 2.635000  0.775000 2.805000 ;
        RECT  1.065000 2.635000  1.235000 2.805000 ;
        RECT  1.525000 2.635000  1.695000 2.805000 ;
        RECT  1.985000 2.635000  2.155000 2.805000 ;
        RECT  2.445000 2.635000  2.615000 2.805000 ;
        RECT  2.905000 2.635000  3.075000 2.805000 ;
        RECT  3.365000 2.635000  3.535000 2.805000 ;
        RECT  3.825000 2.635000  3.995000 2.805000 ;
        RECT  4.285000 2.635000  4.455000 2.805000 ;
        RECT  4.745000 2.635000  4.915000 2.805000 ;
        RECT  5.205000 2.635000  5.375000 2.805000 ;
        RECT  5.665000 2.635000  5.835000 2.805000 ;
        RECT  6.125000 2.635000  6.295000 2.805000 ;
        RECT  6.585000 2.635000  6.755000 2.805000 ;
        RECT  7.045000 2.635000  7.215000 2.805000 ;
        RECT  7.505000 2.635000  7.675000 2.805000 ;
        RECT  7.965000 2.635000  8.135000 2.805000 ;
        RECT  8.425000 2.635000  8.595000 2.805000 ;
        RECT  8.885000 2.635000  9.055000 2.805000 ;
        RECT  9.345000 2.635000  9.515000 2.805000 ;
        RECT  9.805000 2.635000  9.975000 2.805000 ;
        RECT 10.265000 2.635000 10.435000 2.805000 ;
      LAYER met1 ;
        RECT 0.000000 2.480000 10.580000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.090000 0.345000  0.345000 0.635000 ;
      RECT 0.090000 0.635000  0.840000 0.805000 ;
      RECT 0.090000 1.795000  0.840000 1.965000 ;
      RECT 0.090000 1.965000  0.345000 2.465000 ;
      RECT 0.610000 0.805000  0.840000 1.795000 ;
      RECT 1.015000 0.345000  1.185000 2.465000 ;
      RECT 2.045000 0.305000  2.540000 0.475000 ;
      RECT 2.045000 0.475000  2.215000 1.835000 ;
      RECT 2.045000 1.835000  2.440000 2.005000 ;
      RECT 2.270000 2.005000  2.440000 2.135000 ;
      RECT 2.270000 2.135000  2.520000 2.465000 ;
      RECT 2.385000 0.765000  2.735000 1.385000 ;
      RECT 2.610000 1.575000  3.075000 1.965000 ;
      RECT 2.735000 2.135000  3.415000 2.465000 ;
      RECT 2.745000 0.305000  3.600000 0.475000 ;
      RECT 2.905000 0.765000  3.260000 0.985000 ;
      RECT 2.905000 0.985000  3.075000 1.575000 ;
      RECT 3.245000 1.185000  4.935000 1.355000 ;
      RECT 3.245000 1.355000  3.415000 2.135000 ;
      RECT 3.430000 0.475000  3.600000 1.185000 ;
      RECT 3.585000 1.865000  4.660000 2.035000 ;
      RECT 3.585000 2.035000  3.755000 2.375000 ;
      RECT 3.775000 1.525000  5.275000 1.695000 ;
      RECT 4.490000 2.035000  4.660000 2.375000 ;
      RECT 4.765000 1.005000  4.935000 1.185000 ;
      RECT 5.015000 0.275000  5.365000 0.445000 ;
      RECT 5.015000 0.445000  5.275000 0.835000 ;
      RECT 5.105000 0.835000  5.275000 1.525000 ;
      RECT 5.105000 1.695000  5.275000 1.835000 ;
      RECT 5.105000 1.835000  5.665000 2.005000 ;
      RECT 5.465000 0.705000  5.675000 1.495000 ;
      RECT 5.465000 1.495000  6.140000 1.655000 ;
      RECT 5.465000 1.655000  6.430000 1.665000 ;
      RECT 5.495000 2.005000  5.665000 2.465000 ;
      RECT 5.585000 0.255000  6.535000 0.535000 ;
      RECT 5.845000 0.705000  6.195000 1.325000 ;
      RECT 5.900000 2.125000  6.770000 2.465000 ;
      RECT 5.970000 1.665000  6.430000 1.955000 ;
      RECT 6.365000 0.535000  6.535000 1.315000 ;
      RECT 6.365000 1.315000  6.770000 1.485000 ;
      RECT 6.600000 1.485000  6.770000 1.575000 ;
      RECT 6.600000 1.575000  7.820000 1.745000 ;
      RECT 6.600000 1.745000  6.770000 2.125000 ;
      RECT 6.705000 0.695000  7.235000 0.865000 ;
      RECT 6.705000 0.865000  6.925000 1.145000 ;
      RECT 7.065000 0.295000  8.135000 0.465000 ;
      RECT 7.065000 0.465000  7.235000 0.695000 ;
      RECT 7.360000 1.915000  8.160000 2.085000 ;
      RECT 7.360000 2.085000  7.530000 2.375000 ;
      RECT 7.815000 0.465000  8.135000 0.820000 ;
      RECT 7.815000 0.820000  8.140000 0.995000 ;
      RECT 7.815000 0.995000  8.435000 1.295000 ;
      RECT 7.990000 1.295000  8.435000 1.325000 ;
      RECT 7.990000 1.325000  8.160000 1.915000 ;
      RECT 9.195000 0.345000  9.445000 0.995000 ;
      RECT 9.195000 0.995000 10.055000 1.325000 ;
      RECT 9.195000 1.325000  9.525000 2.425000 ;
    LAYER mcon ;
      RECT 0.610000 1.105000 0.780000 1.275000 ;
      RECT 1.015000 1.785000 1.185000 1.955000 ;
      RECT 2.445000 1.105000 2.615000 1.275000 ;
      RECT 2.905000 1.785000 3.075000 1.955000 ;
      RECT 6.025000 1.105000 6.195000 1.275000 ;
      RECT 6.025000 1.785000 6.195000 1.955000 ;
    LAYER met1 ;
      RECT 0.550000 1.075000 0.840000 1.120000 ;
      RECT 0.550000 1.120000 6.255000 1.260000 ;
      RECT 0.550000 1.260000 0.840000 1.305000 ;
      RECT 0.955000 1.755000 1.245000 1.800000 ;
      RECT 0.955000 1.800000 6.255000 1.940000 ;
      RECT 0.955000 1.940000 1.245000 1.985000 ;
      RECT 2.385000 1.075000 2.675000 1.120000 ;
      RECT 2.385000 1.260000 2.675000 1.305000 ;
      RECT 2.845000 1.755000 3.135000 1.800000 ;
      RECT 2.845000 1.940000 3.135000 1.985000 ;
      RECT 5.965000 1.075000 6.255000 1.120000 ;
      RECT 5.965000 1.260000 6.255000 1.305000 ;
      RECT 5.965000 1.755000 6.255000 1.800000 ;
      RECT 5.965000 1.940000 6.255000 1.985000 ;
  END
END sky130_fd_sc_hd__dfrbp_1
END LIBRARY
