# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hd__lpflow_clkinvkapwr_8
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_hd__lpflow_clkinvkapwr_8 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  5.980000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  2.304000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.455000 1.035000 4.865000 1.290000 ;
    END
  END A
  PIN Y
    ANTENNADIFFAREA  2.090400 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.115000 0.695000 5.440000 0.865000 ;
        RECT 0.115000 0.865000 0.285000 1.460000 ;
        RECT 0.115000 1.460000 5.440000 1.630000 ;
        RECT 0.595000 1.630000 0.765000 2.435000 ;
        RECT 1.440000 1.630000 1.610000 2.435000 ;
        RECT 1.535000 0.280000 1.725000 0.695000 ;
        RECT 2.280000 1.630000 2.450000 2.435000 ;
        RECT 2.395000 0.280000 2.585000 0.695000 ;
        RECT 3.120000 1.630000 3.290000 2.435000 ;
        RECT 3.255000 0.280000 3.445000 0.695000 ;
        RECT 3.960000 1.630000 4.130000 2.435000 ;
        RECT 4.115000 0.280000 4.305000 0.695000 ;
        RECT 4.800000 1.630000 4.970000 2.435000 ;
        RECT 5.170000 0.865000 5.440000 1.460000 ;
    END
  END Y
  PIN KAPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.095000 1.800000 0.425000 2.465000 ;
        RECT 0.940000 1.800000 1.270000 2.465000 ;
        RECT 1.780000 1.800000 2.110000 2.465000 ;
        RECT 2.620000 1.800000 2.950000 2.465000 ;
        RECT 3.460000 1.800000 3.790000 2.465000 ;
        RECT 4.300000 1.800000 4.630000 2.465000 ;
        RECT 5.140000 1.800000 5.470000 2.465000 ;
      LAYER mcon ;
        RECT 0.130000 2.125000 0.300000 2.295000 ;
        RECT 0.990000 2.125000 1.160000 2.295000 ;
        RECT 1.890000 2.125000 2.060000 2.295000 ;
        RECT 2.770000 2.125000 2.940000 2.295000 ;
        RECT 3.495000 2.125000 3.665000 2.295000 ;
        RECT 4.355000 2.125000 4.525000 2.295000 ;
        RECT 5.255000 2.125000 5.425000 2.295000 ;
      LAYER met1 ;
        RECT 0.070000 2.080000 0.360000 2.140000 ;
        RECT 0.070000 2.140000 5.910000 2.340000 ;
        RECT 0.930000 2.080000 1.220000 2.140000 ;
        RECT 1.830000 2.080000 2.120000 2.140000 ;
        RECT 2.710000 2.080000 3.000000 2.140000 ;
        RECT 3.435000 2.080000 3.725000 2.140000 ;
        RECT 4.295000 2.080000 4.585000 2.140000 ;
        RECT 5.195000 2.080000 5.485000 2.140000 ;
    END
  END KAPWR
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 5.980000 0.085000 ;
        RECT 1.035000  0.085000 1.365000 0.525000 ;
        RECT 1.895000  0.085000 2.225000 0.525000 ;
        RECT 2.755000  0.085000 3.085000 0.525000 ;
        RECT 3.615000  0.085000 3.945000 0.525000 ;
        RECT 4.475000  0.085000 4.805000 0.525000 ;
      LAYER mcon ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
        RECT 0.605000 -0.085000 0.775000 0.085000 ;
        RECT 1.065000 -0.085000 1.235000 0.085000 ;
        RECT 1.525000 -0.085000 1.695000 0.085000 ;
        RECT 1.985000 -0.085000 2.155000 0.085000 ;
        RECT 2.445000 -0.085000 2.615000 0.085000 ;
        RECT 2.905000 -0.085000 3.075000 0.085000 ;
        RECT 3.365000 -0.085000 3.535000 0.085000 ;
        RECT 3.825000 -0.085000 3.995000 0.085000 ;
        RECT 4.285000 -0.085000 4.455000 0.085000 ;
        RECT 4.745000 -0.085000 4.915000 0.085000 ;
        RECT 5.205000 -0.085000 5.375000 0.085000 ;
        RECT 5.665000 -0.085000 5.835000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.240000 5.980000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 5.980000 2.805000 ;
      LAYER mcon ;
        RECT 0.145000 2.635000 0.315000 2.805000 ;
        RECT 0.605000 2.635000 0.775000 2.805000 ;
        RECT 1.065000 2.635000 1.235000 2.805000 ;
        RECT 1.525000 2.635000 1.695000 2.805000 ;
        RECT 1.985000 2.635000 2.155000 2.805000 ;
        RECT 2.445000 2.635000 2.615000 2.805000 ;
        RECT 2.905000 2.635000 3.075000 2.805000 ;
        RECT 3.365000 2.635000 3.535000 2.805000 ;
        RECT 3.825000 2.635000 3.995000 2.805000 ;
        RECT 4.285000 2.635000 4.455000 2.805000 ;
        RECT 4.745000 2.635000 4.915000 2.805000 ;
        RECT 5.205000 2.635000 5.375000 2.805000 ;
        RECT 5.665000 2.635000 5.835000 2.805000 ;
      LAYER met1 ;
        RECT 0.000000 2.480000 5.980000 2.960000 ;
    END
  END VPWR
END sky130_fd_sc_hd__lpflow_clkinvkapwr_8
END LIBRARY
