# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hd__edfxtp_1
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_hd__edfxtp_1 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  11.04000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN D
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.695000 0.765000 1.915000 1.720000 ;
    END
  END D
  PIN DE
    ANTENNAGATEAREA  0.318000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.110000 0.765000 2.565000 1.185000 ;
        RECT 2.110000 1.185000 2.325000 1.370000 ;
    END
  END DE
  PIN Q
    ANTENNADIFFAREA  0.462000 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 10.465000 0.305000 10.795000 2.420000 ;
    END
  END Q
  PIN CLK
    ANTENNAGATEAREA  0.159000 ;
    DIRECTION INPUT ;
    USE CLOCK ;
    PORT
      LAYER li1 ;
        RECT 0.095000 0.975000 0.445000 1.625000 ;
    END
  END CLK
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT  0.000000 -0.085000 11.040000 0.085000 ;
        RECT  0.515000  0.085000  0.845000 0.465000 ;
        RECT  2.235000  0.085000  2.565000 0.515000 ;
        RECT  3.185000  0.085000  3.515000 0.610000 ;
        RECT  5.945000  0.085000  6.340000 0.560000 ;
        RECT  7.165000  0.085000  7.440000 0.615000 ;
        RECT  9.050000  0.085000  9.365000 0.615000 ;
        RECT 10.050000  0.085000 10.295000 0.900000 ;
      LAYER mcon ;
        RECT  0.145000 -0.085000  0.315000 0.085000 ;
        RECT  0.605000 -0.085000  0.775000 0.085000 ;
        RECT  1.065000 -0.085000  1.235000 0.085000 ;
        RECT  1.525000 -0.085000  1.695000 0.085000 ;
        RECT  1.985000 -0.085000  2.155000 0.085000 ;
        RECT  2.445000 -0.085000  2.615000 0.085000 ;
        RECT  2.905000 -0.085000  3.075000 0.085000 ;
        RECT  3.365000 -0.085000  3.535000 0.085000 ;
        RECT  3.825000 -0.085000  3.995000 0.085000 ;
        RECT  4.285000 -0.085000  4.455000 0.085000 ;
        RECT  4.745000 -0.085000  4.915000 0.085000 ;
        RECT  5.205000 -0.085000  5.375000 0.085000 ;
        RECT  5.665000 -0.085000  5.835000 0.085000 ;
        RECT  6.125000 -0.085000  6.295000 0.085000 ;
        RECT  6.585000 -0.085000  6.755000 0.085000 ;
        RECT  7.045000 -0.085000  7.215000 0.085000 ;
        RECT  7.505000 -0.085000  7.675000 0.085000 ;
        RECT  7.965000 -0.085000  8.135000 0.085000 ;
        RECT  8.425000 -0.085000  8.595000 0.085000 ;
        RECT  8.885000 -0.085000  9.055000 0.085000 ;
        RECT  9.345000 -0.085000  9.515000 0.085000 ;
        RECT  9.805000 -0.085000  9.975000 0.085000 ;
        RECT 10.265000 -0.085000 10.435000 0.085000 ;
        RECT 10.725000 -0.085000 10.895000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.240000 11.040000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT  0.000000 2.635000 11.040000 2.805000 ;
        RECT  0.515000 2.135000  0.845000 2.635000 ;
        RECT  2.235000 1.890000  2.565000 2.635000 ;
        RECT  3.265000 1.825000  3.460000 2.635000 ;
        RECT  6.125000 1.835000  6.360000 2.635000 ;
        RECT  7.070000 2.105000  7.360000 2.635000 ;
        RECT  8.980000 2.135000  9.240000 2.635000 ;
        RECT 10.050000 1.465000 10.295000 2.635000 ;
      LAYER mcon ;
        RECT  0.145000 2.635000  0.315000 2.805000 ;
        RECT  0.605000 2.635000  0.775000 2.805000 ;
        RECT  1.065000 2.635000  1.235000 2.805000 ;
        RECT  1.525000 2.635000  1.695000 2.805000 ;
        RECT  1.985000 2.635000  2.155000 2.805000 ;
        RECT  2.445000 2.635000  2.615000 2.805000 ;
        RECT  2.905000 2.635000  3.075000 2.805000 ;
        RECT  3.365000 2.635000  3.535000 2.805000 ;
        RECT  3.825000 2.635000  3.995000 2.805000 ;
        RECT  4.285000 2.635000  4.455000 2.805000 ;
        RECT  4.745000 2.635000  4.915000 2.805000 ;
        RECT  5.205000 2.635000  5.375000 2.805000 ;
        RECT  5.665000 2.635000  5.835000 2.805000 ;
        RECT  6.125000 2.635000  6.295000 2.805000 ;
        RECT  6.585000 2.635000  6.755000 2.805000 ;
        RECT  7.045000 2.635000  7.215000 2.805000 ;
        RECT  7.505000 2.635000  7.675000 2.805000 ;
        RECT  7.965000 2.635000  8.135000 2.805000 ;
        RECT  8.425000 2.635000  8.595000 2.805000 ;
        RECT  8.885000 2.635000  9.055000 2.805000 ;
        RECT  9.345000 2.635000  9.515000 2.805000 ;
        RECT  9.805000 2.635000  9.975000 2.805000 ;
        RECT 10.265000 2.635000 10.435000 2.805000 ;
        RECT 10.725000 2.635000 10.895000 2.805000 ;
      LAYER met1 ;
        RECT 0.000000 2.480000 11.040000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.175000 0.345000 0.345000 0.635000 ;
      RECT 0.175000 0.635000 0.845000 0.805000 ;
      RECT 0.175000 1.795000 0.845000 1.965000 ;
      RECT 0.175000 1.965000 0.345000 2.465000 ;
      RECT 0.615000 0.805000 0.845000 1.795000 ;
      RECT 1.015000 0.345000 1.185000 2.465000 ;
      RECT 1.355000 0.255000 1.785000 0.515000 ;
      RECT 1.355000 0.515000 1.525000 1.890000 ;
      RECT 1.355000 1.890000 1.785000 2.465000 ;
      RECT 2.495000 1.355000 3.085000 1.720000 ;
      RECT 2.755000 1.720000 3.085000 2.425000 ;
      RECT 2.780000 0.255000 3.005000 0.845000 ;
      RECT 2.780000 0.845000 3.635000 1.175000 ;
      RECT 2.780000 1.175000 3.085000 1.355000 ;
      RECT 3.805000 0.685000 3.975000 1.320000 ;
      RECT 3.805000 1.320000 4.175000 1.650000 ;
      RECT 4.125000 1.820000 4.515000 2.020000 ;
      RECT 4.125000 2.020000 4.455000 2.465000 ;
      RECT 4.145000 0.255000 4.415000 0.980000 ;
      RECT 4.145000 0.980000 4.515000 1.150000 ;
      RECT 4.345000 1.150000 4.515000 1.820000 ;
      RECT 4.795000 1.125000 4.980000 1.720000 ;
      RECT 4.815000 0.735000 5.320000 0.955000 ;
      RECT 4.915000 2.175000 5.955000 2.375000 ;
      RECT 5.005000 0.255000 5.680000 0.565000 ;
      RECT 5.150000 0.955000 5.320000 1.655000 ;
      RECT 5.150000 1.655000 5.615000 2.005000 ;
      RECT 5.510000 0.565000 5.680000 1.315000 ;
      RECT 5.510000 1.315000 6.360000 1.485000 ;
      RECT 5.785000 1.485000 6.360000 1.575000 ;
      RECT 5.785000 1.575000 5.955000 2.175000 ;
      RECT 5.870000 0.765000 6.935000 1.045000 ;
      RECT 5.870000 1.045000 7.445000 1.065000 ;
      RECT 5.870000 1.065000 6.070000 1.095000 ;
      RECT 6.190000 1.245000 6.360000 1.315000 ;
      RECT 6.530000 0.255000 6.935000 0.765000 ;
      RECT 6.530000 1.065000 7.445000 1.375000 ;
      RECT 6.530000 1.375000 6.860000 2.465000 ;
      RECT 7.790000 1.245000 7.980000 1.965000 ;
      RECT 7.925000 2.165000 8.810000 2.355000 ;
      RECT 8.005000 0.705000 8.470000 1.035000 ;
      RECT 8.025000 0.330000 8.810000 0.535000 ;
      RECT 8.150000 1.035000 8.470000 1.995000 ;
      RECT 8.640000 0.535000 8.810000 0.995000 ;
      RECT 8.640000 0.995000 9.510000 1.325000 ;
      RECT 8.640000 1.325000 8.810000 2.165000 ;
      RECT 8.980000 1.530000 9.880000 1.905000 ;
      RECT 9.540000 1.905000 9.880000 2.465000 ;
      RECT 9.550000 0.300000 9.880000 0.825000 ;
      RECT 9.690000 0.825000 9.880000 1.530000 ;
    LAYER mcon ;
      RECT 0.635000 1.785000 0.805000 1.955000 ;
      RECT 1.015000 1.445000 1.185000 1.615000 ;
      RECT 1.355000 0.425000 1.525000 0.595000 ;
      RECT 3.805000 0.765000 3.975000 0.935000 ;
      RECT 4.185000 0.425000 4.355000 0.595000 ;
      RECT 4.800000 1.445000 4.970000 1.615000 ;
      RECT 5.210000 1.785000 5.380000 1.955000 ;
      RECT 7.800000 1.785000 7.970000 1.955000 ;
      RECT 8.220000 1.445000 8.390000 1.615000 ;
      RECT 9.700000 0.765000 9.870000 0.935000 ;
    LAYER met1 ;
      RECT 0.575000 1.755000 0.865000 1.800000 ;
      RECT 0.575000 1.800000 8.030000 1.940000 ;
      RECT 0.575000 1.940000 0.865000 1.985000 ;
      RECT 0.955000 1.415000 1.245000 1.460000 ;
      RECT 0.955000 1.460000 8.450000 1.600000 ;
      RECT 0.955000 1.600000 1.245000 1.645000 ;
      RECT 1.295000 0.395000 4.415000 0.580000 ;
      RECT 1.295000 0.580000 1.585000 0.625000 ;
      RECT 3.745000 0.735000 4.035000 0.780000 ;
      RECT 3.745000 0.780000 9.930000 0.920000 ;
      RECT 3.745000 0.920000 4.035000 0.965000 ;
      RECT 4.125000 0.580000 4.415000 0.625000 ;
      RECT 4.740000 1.415000 5.030000 1.460000 ;
      RECT 4.740000 1.600000 5.030000 1.645000 ;
      RECT 5.150000 1.755000 5.440000 1.800000 ;
      RECT 5.150000 1.940000 5.440000 1.985000 ;
      RECT 7.740000 1.755000 8.030000 1.800000 ;
      RECT 7.740000 1.940000 8.030000 1.985000 ;
      RECT 8.160000 1.415000 8.450000 1.460000 ;
      RECT 8.160000 1.600000 8.450000 1.645000 ;
      RECT 9.640000 0.735000 9.930000 0.780000 ;
      RECT 9.640000 0.920000 9.930000 0.965000 ;
  END
END sky130_fd_sc_hd__edfxtp_1
END LIBRARY
