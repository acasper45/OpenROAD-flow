# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hd__xor3_2
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_hd__xor3_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  9.200000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.246000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.965000 1.075000 8.375000 1.325000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.661500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 7.145000 0.995000 7.315000 1.445000 ;
        RECT 7.145000 1.445000 7.725000 1.615000 ;
    END
  END B
  PIN C
    ANTENNAGATEAREA  0.381000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 2.320000 0.995000 2.955000 1.325000 ;
    END
  END C
  PIN X
    ANTENNADIFFAREA  0.445500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.545000 0.660000 1.050000 0.925000 ;
        RECT 0.545000 0.925000 0.860000 1.440000 ;
        RECT 0.545000 1.440000 1.070000 2.045000 ;
        RECT 0.800000 0.350000 1.050000 0.660000 ;
        RECT 0.820000 2.045000 1.070000 2.465000 ;
    END
  END X
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 9.200000 0.085000 ;
        RECT 0.300000  0.085000 0.630000 0.465000 ;
        RECT 1.220000  0.085000 1.470000 0.525000 ;
        RECT 4.390000  0.085000 4.560000 0.865000 ;
        RECT 8.395000  0.085000 8.565000 0.565000 ;
      LAYER mcon ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
        RECT 0.605000 -0.085000 0.775000 0.085000 ;
        RECT 1.065000 -0.085000 1.235000 0.085000 ;
        RECT 1.525000 -0.085000 1.695000 0.085000 ;
        RECT 1.985000 -0.085000 2.155000 0.085000 ;
        RECT 2.445000 -0.085000 2.615000 0.085000 ;
        RECT 2.905000 -0.085000 3.075000 0.085000 ;
        RECT 3.365000 -0.085000 3.535000 0.085000 ;
        RECT 3.825000 -0.085000 3.995000 0.085000 ;
        RECT 4.285000 -0.085000 4.455000 0.085000 ;
        RECT 4.745000 -0.085000 4.915000 0.085000 ;
        RECT 5.205000 -0.085000 5.375000 0.085000 ;
        RECT 5.665000 -0.085000 5.835000 0.085000 ;
        RECT 6.125000 -0.085000 6.295000 0.085000 ;
        RECT 6.585000 -0.085000 6.755000 0.085000 ;
        RECT 7.045000 -0.085000 7.215000 0.085000 ;
        RECT 7.505000 -0.085000 7.675000 0.085000 ;
        RECT 7.965000 -0.085000 8.135000 0.085000 ;
        RECT 8.425000 -0.085000 8.595000 0.085000 ;
        RECT 8.885000 -0.085000 9.055000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.240000 9.200000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 9.200000 2.805000 ;
        RECT 0.300000 2.215000 0.650000 2.635000 ;
        RECT 1.240000 2.215000 1.575000 2.635000 ;
        RECT 4.145000 2.235000 4.475000 2.635000 ;
        RECT 8.315000 2.275000 8.650000 2.635000 ;
      LAYER mcon ;
        RECT 0.145000 2.635000 0.315000 2.805000 ;
        RECT 0.605000 2.635000 0.775000 2.805000 ;
        RECT 1.065000 2.635000 1.235000 2.805000 ;
        RECT 1.525000 2.635000 1.695000 2.805000 ;
        RECT 1.985000 2.635000 2.155000 2.805000 ;
        RECT 2.445000 2.635000 2.615000 2.805000 ;
        RECT 2.905000 2.635000 3.075000 2.805000 ;
        RECT 3.365000 2.635000 3.535000 2.805000 ;
        RECT 3.825000 2.635000 3.995000 2.805000 ;
        RECT 4.285000 2.635000 4.455000 2.805000 ;
        RECT 4.745000 2.635000 4.915000 2.805000 ;
        RECT 5.205000 2.635000 5.375000 2.805000 ;
        RECT 5.665000 2.635000 5.835000 2.805000 ;
        RECT 6.125000 2.635000 6.295000 2.805000 ;
        RECT 6.585000 2.635000 6.755000 2.805000 ;
        RECT 7.045000 2.635000 7.215000 2.805000 ;
        RECT 7.505000 2.635000 7.675000 2.805000 ;
        RECT 7.965000 2.635000 8.135000 2.805000 ;
        RECT 8.425000 2.635000 8.595000 2.805000 ;
        RECT 8.885000 2.635000 9.055000 2.805000 ;
      LAYER met1 ;
        RECT 0.000000 2.480000 9.200000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 1.210000 0.995000 1.410000 1.325000 ;
      RECT 1.240000 0.695000 1.810000 0.865000 ;
      RECT 1.240000 0.865000 1.410000 0.995000 ;
      RECT 1.240000 1.325000 1.410000 1.875000 ;
      RECT 1.240000 1.875000 1.930000 2.045000 ;
      RECT 1.640000 0.255000 3.200000 0.425000 ;
      RECT 1.640000 0.425000 1.810000 0.695000 ;
      RECT 1.645000 1.535000 3.295000 1.705000 ;
      RECT 1.760000 2.045000 1.930000 2.235000 ;
      RECT 1.760000 2.235000 3.355000 2.405000 ;
      RECT 1.980000 0.595000 2.150000 1.535000 ;
      RECT 2.330000 1.895000 3.635000 2.065000 ;
      RECT 2.430000 0.655000 3.540000 0.825000 ;
      RECT 2.850000 0.425000 3.200000 0.455000 ;
      RECT 3.125000 0.995000 3.400000 1.325000 ;
      RECT 3.125000 1.325000 3.295000 1.535000 ;
      RECT 3.370000 0.255000 4.220000 0.425000 ;
      RECT 3.370000 0.425000 3.540000 0.655000 ;
      RECT 3.465000 1.525000 3.995000 1.695000 ;
      RECT 3.465000 1.695000 3.635000 1.895000 ;
      RECT 3.570000 2.235000 3.975000 2.405000 ;
      RECT 3.710000 0.595000 3.880000 1.375000 ;
      RECT 3.710000 1.375000 3.995000 1.525000 ;
      RECT 3.805000 1.895000 4.980000 2.065000 ;
      RECT 3.805000 2.065000 3.975000 2.235000 ;
      RECT 4.050000 0.425000 4.220000 1.035000 ;
      RECT 4.050000 1.035000 4.335000 1.205000 ;
      RECT 4.165000 1.205000 4.335000 1.895000 ;
      RECT 4.565000 1.445000 4.980000 1.715000 ;
      RECT 4.740000 0.415000 4.980000 1.445000 ;
      RECT 4.810000 2.065000 4.980000 2.275000 ;
      RECT 4.810000 2.275000 7.905000 2.445000 ;
      RECT 5.155000 0.265000 5.570000 0.485000 ;
      RECT 5.155000 0.485000 5.375000 0.595000 ;
      RECT 5.155000 0.595000 5.325000 2.105000 ;
      RECT 5.495000 0.720000 5.910000 0.825000 ;
      RECT 5.495000 0.825000 5.715000 0.890000 ;
      RECT 5.495000 0.890000 5.665000 2.275000 ;
      RECT 5.545000 0.655000 5.910000 0.720000 ;
      RECT 5.740000 0.320000 5.910000 0.655000 ;
      RECT 5.855000 1.445000 6.635000 1.615000 ;
      RECT 5.855000 1.615000 6.270000 2.045000 ;
      RECT 5.870000 0.995000 6.295000 1.270000 ;
      RECT 6.080000 0.630000 6.295000 0.995000 ;
      RECT 6.465000 0.255000 7.610000 0.425000 ;
      RECT 6.465000 0.425000 6.635000 1.445000 ;
      RECT 6.805000 0.595000 6.975000 1.935000 ;
      RECT 6.805000 1.935000 9.115000 2.105000 ;
      RECT 7.145000 0.425000 7.610000 0.465000 ;
      RECT 7.485000 0.730000 7.690000 0.945000 ;
      RECT 7.485000 0.945000 7.795000 1.275000 ;
      RECT 7.895000 1.495000 8.715000 1.705000 ;
      RECT 7.935000 0.295000 8.225000 0.735000 ;
      RECT 7.935000 0.735000 8.715000 0.750000 ;
      RECT 7.975000 0.750000 8.715000 0.905000 ;
      RECT 8.545000 0.905000 8.715000 0.995000 ;
      RECT 8.545000 0.995000 8.775000 1.325000 ;
      RECT 8.545000 1.325000 8.715000 1.495000 ;
      RECT 8.630000 1.875000 9.115000 1.935000 ;
      RECT 8.815000 0.255000 9.115000 0.585000 ;
      RECT 8.820000 2.105000 9.115000 2.465000 ;
      RECT 8.945000 0.585000 9.115000 1.875000 ;
    LAYER mcon ;
      RECT 3.825000 1.445000 3.995000 1.615000 ;
      RECT 4.745000 0.765000 4.915000 0.935000 ;
      RECT 5.205000 0.425000 5.375000 0.595000 ;
      RECT 6.125000 0.765000 6.295000 0.935000 ;
      RECT 6.125000 1.445000 6.295000 1.615000 ;
      RECT 7.505000 0.765000 7.675000 0.935000 ;
      RECT 7.965000 0.425000 8.135000 0.595000 ;
    LAYER met1 ;
      RECT 3.765000 1.415000 4.055000 1.460000 ;
      RECT 3.765000 1.460000 6.355000 1.600000 ;
      RECT 3.765000 1.600000 4.055000 1.645000 ;
      RECT 4.685000 0.735000 4.975000 0.780000 ;
      RECT 4.685000 0.780000 7.735000 0.920000 ;
      RECT 4.685000 0.920000 4.975000 0.965000 ;
      RECT 5.145000 0.395000 5.435000 0.440000 ;
      RECT 5.145000 0.440000 8.195000 0.580000 ;
      RECT 5.145000 0.580000 5.435000 0.625000 ;
      RECT 6.065000 0.735000 6.355000 0.780000 ;
      RECT 6.065000 0.920000 6.355000 0.965000 ;
      RECT 6.065000 1.415000 6.355000 1.460000 ;
      RECT 6.065000 1.600000 6.355000 1.645000 ;
      RECT 7.445000 0.735000 7.735000 0.780000 ;
      RECT 7.445000 0.920000 7.735000 0.965000 ;
      RECT 7.905000 0.395000 8.195000 0.440000 ;
      RECT 7.905000 0.580000 8.195000 0.625000 ;
  END
END sky130_fd_sc_hd__xor3_2
END LIBRARY
