# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hd__nor3b_2
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_hd__nor3b_2 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  4.600000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.110000 1.075000 0.965000 1.285000 ;
    END
  END A
  PIN B
    ANTENNAGATEAREA  0.495000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 1.135000 1.075000 2.640000 1.285000 ;
    END
  END B
  PIN C_N
    ANTENNAGATEAREA  0.126000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 4.030000 1.075000 4.515000 1.285000 ;
    END
  END C_N
  PIN Y
    ANTENNADIFFAREA  0.796500 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.535000 0.255000 0.865000 0.725000 ;
        RECT 0.535000 0.725000 3.105000 0.905000 ;
        RECT 1.375000 0.255000 1.705000 0.725000 ;
        RECT 2.775000 0.255000 3.105000 0.725000 ;
        RECT 2.815000 0.905000 3.065000 2.125000 ;
    END
  END Y
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT 0.000000 -0.085000 4.600000 0.085000 ;
        RECT 0.090000  0.085000 0.365000 0.905000 ;
        RECT 1.035000  0.085000 1.205000 0.555000 ;
        RECT 1.875000  0.085000 2.605000 0.555000 ;
        RECT 3.275000  0.085000 3.480000 0.895000 ;
        RECT 4.215000  0.085000 4.505000 0.825000 ;
      LAYER mcon ;
        RECT 0.145000 -0.085000 0.315000 0.085000 ;
        RECT 0.605000 -0.085000 0.775000 0.085000 ;
        RECT 1.065000 -0.085000 1.235000 0.085000 ;
        RECT 1.525000 -0.085000 1.695000 0.085000 ;
        RECT 1.985000 -0.085000 2.155000 0.085000 ;
        RECT 2.445000 -0.085000 2.615000 0.085000 ;
        RECT 2.905000 -0.085000 3.075000 0.085000 ;
        RECT 3.365000 -0.085000 3.535000 0.085000 ;
        RECT 3.825000 -0.085000 3.995000 0.085000 ;
        RECT 4.285000 -0.085000 4.455000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.240000 4.600000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 4.600000 2.805000 ;
        RECT 0.575000 1.795000 0.825000 2.635000 ;
        RECT 4.215000 1.540000 4.465000 2.635000 ;
      LAYER mcon ;
        RECT 0.145000 2.635000 0.315000 2.805000 ;
        RECT 0.605000 2.635000 0.775000 2.805000 ;
        RECT 1.065000 2.635000 1.235000 2.805000 ;
        RECT 1.525000 2.635000 1.695000 2.805000 ;
        RECT 1.985000 2.635000 2.155000 2.805000 ;
        RECT 2.445000 2.635000 2.615000 2.805000 ;
        RECT 2.905000 2.635000 3.075000 2.805000 ;
        RECT 3.365000 2.635000 3.535000 2.805000 ;
        RECT 3.825000 2.635000 3.995000 2.805000 ;
        RECT 4.285000 2.635000 4.455000 2.805000 ;
      LAYER met1 ;
        RECT 0.000000 2.480000 4.600000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.090000 1.455000 2.085000 1.625000 ;
      RECT 0.090000 1.625000 0.405000 2.465000 ;
      RECT 0.995000 1.625000 1.245000 2.465000 ;
      RECT 1.415000 1.795000 1.665000 2.295000 ;
      RECT 1.415000 2.295000 3.480000 2.465000 ;
      RECT 1.835000 1.625000 2.085000 2.125000 ;
      RECT 2.375000 1.455000 2.645000 2.295000 ;
      RECT 3.235000 1.075000 3.860000 1.285000 ;
      RECT 3.235000 1.455000 3.480000 2.295000 ;
      RECT 3.690000 0.380000 4.045000 0.905000 ;
      RECT 3.690000 0.905000 3.860000 1.075000 ;
      RECT 3.690000 1.285000 3.860000 1.455000 ;
      RECT 3.690000 1.455000 4.045000 1.870000 ;
  END
END sky130_fd_sc_hd__nor3b_2
END LIBRARY
