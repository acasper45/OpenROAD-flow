# Copyright 2020 The SkyWater PDK Authors
#
# Licensed under the Apache License, Version 2.0 (the "License");
# you may not use this file except in compliance with the License.
# You may obtain a copy of the License at
#
#     https://www.apache.org/licenses/LICENSE-2.0
#
# Unless required by applicable law or agreed to in writing, software
# distributed under the License is distributed on an "AS IS" BASIS,
# WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
# See the License for the specific language governing permissions and
# limitations under the License.
#
# SPDX-License-Identifier: Apache-2.0

VERSION 5.7 ;
  NAMESCASESENSITIVE ON ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
UNITS
  DATABASE MICRONS 200 ;
END UNITS
MACRO sky130_fd_sc_hd__lpflow_isobufsrckapwr_16
  CLASS CORE ;
  SOURCE USER ;
  FOREIGN sky130_fd_sc_hd__lpflow_isobufsrckapwr_16 ;
  ORIGIN  0.000000  0.000000 ;
  SIZE  14.26000 BY  2.720000 ;
  SYMMETRY X Y R90 ;
  SITE unithd ;
  PIN A
    ANTENNAGATEAREA  0.247500 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 0.085000 1.075000 0.615000 1.320000 ;
    END
  END A
  PIN SLEEP
    ANTENNAGATEAREA  0.990000 ;
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT 3.260000 1.075000 4.700000 1.275000 ;
    END
  END SLEEP
  PIN X
    ANTENNADIFFAREA  3.180800 ;
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER li1 ;
        RECT  7.340000 0.280000  7.600000 0.735000 ;
        RECT  7.340000 0.735000 14.085000 0.905000 ;
        RECT  7.375000 1.495000 14.085000 1.720000 ;
        RECT  7.375000 1.720000 12.745000 1.735000 ;
        RECT  7.375000 1.735000  7.600000 2.460000 ;
        RECT  8.200000 0.280000  8.460000 0.735000 ;
        RECT  8.200000 1.735000  8.460000 2.460000 ;
        RECT  9.060000 0.280000  9.320000 0.735000 ;
        RECT  9.060000 1.735000  9.320000 2.460000 ;
        RECT  9.905000 0.280000 10.180000 0.735000 ;
        RECT  9.920000 1.735000 10.180000 2.460000 ;
        RECT 10.765000 0.280000 11.025000 0.735000 ;
        RECT 10.765000 1.735000 11.025000 2.460000 ;
        RECT 11.625000 0.280000 11.885000 0.735000 ;
        RECT 11.625000 1.735000 11.885000 2.460000 ;
        RECT 12.485000 0.280000 12.745000 0.735000 ;
        RECT 12.485000 1.735000 12.745000 2.460000 ;
        RECT 12.920000 0.905000 14.085000 1.495000 ;
        RECT 13.355000 0.280000 13.615000 0.735000 ;
        RECT 13.355000 1.720000 13.645000 2.460000 ;
    END
  END X
  PIN KAPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT  5.155000 1.495000  5.485000 2.465000 ;
        RECT  6.015000 1.495000  6.345000 2.465000 ;
        RECT  6.875000 1.495000  7.205000 2.465000 ;
        RECT  7.770000 1.905000  8.030000 2.465000 ;
        RECT  8.630000 1.905000  8.890000 2.465000 ;
        RECT  9.490000 1.905000  9.750000 2.465000 ;
        RECT 10.350000 1.905000 10.595000 2.465000 ;
        RECT 11.210000 1.905000 11.455000 2.465000 ;
        RECT 12.070000 1.905000 12.315000 2.465000 ;
        RECT 12.930000 1.905000 13.185000 2.465000 ;
        RECT 13.815000 1.890000 14.085000 2.465000 ;
      LAYER mcon ;
        RECT  5.235000 2.125000  5.405000 2.295000 ;
        RECT  6.095000 2.125000  6.265000 2.295000 ;
        RECT  6.950000 2.125000  7.120000 2.295000 ;
        RECT  7.800000 2.125000  7.970000 2.295000 ;
        RECT  8.680000 2.125000  8.850000 2.295000 ;
        RECT  9.540000 2.125000  9.710000 2.295000 ;
        RECT 10.395000 2.125000 10.565000 2.295000 ;
        RECT 11.255000 2.125000 11.425000 2.295000 ;
        RECT 12.110000 2.125000 12.280000 2.295000 ;
        RECT 12.960000 2.125000 13.130000 2.295000 ;
        RECT 13.840000 2.125000 14.010000 2.295000 ;
      LAYER met1 ;
        RECT  0.070000 2.140000 14.190000 2.340000 ;
        RECT  5.175000 2.080000  5.465000 2.140000 ;
        RECT  6.035000 2.080000  6.325000 2.140000 ;
        RECT  6.890000 2.080000  7.180000 2.140000 ;
        RECT  7.740000 2.080000  8.030000 2.140000 ;
        RECT  8.620000 2.080000  8.910000 2.140000 ;
        RECT  9.480000 2.080000  9.770000 2.140000 ;
        RECT 10.335000 2.080000 10.625000 2.140000 ;
        RECT 11.195000 2.080000 11.485000 2.140000 ;
        RECT 12.050000 2.080000 12.340000 2.140000 ;
        RECT 12.900000 2.080000 13.190000 2.140000 ;
        RECT 13.780000 2.080000 14.070000 2.140000 ;
    END
  END KAPWR
  PIN VGND
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE GROUND ;
    PORT
      LAYER li1 ;
        RECT  0.000000 -0.085000 14.260000 0.085000 ;
        RECT  0.245000  0.085000  0.535000 0.905000 ;
        RECT  1.215000  0.085000  1.505000 0.905000 ;
        RECT  2.175000  0.085000  2.345000 0.555000 ;
        RECT  3.015000  0.085000  3.185000 0.555000 ;
        RECT  3.855000  0.085000  4.025000 0.555000 ;
        RECT  4.695000  0.085000  5.450000 0.565000 ;
        RECT  4.695000  0.565000  4.975000 0.905000 ;
        RECT  6.050000  0.085000  6.310000 0.610000 ;
        RECT  6.910000  0.085000  7.170000 0.645000 ;
        RECT  7.770000  0.085000  8.030000 0.565000 ;
        RECT  8.630000  0.085000  8.890000 0.565000 ;
        RECT  9.490000  0.085000  9.735000 0.565000 ;
        RECT 10.350000  0.085000 10.595000 0.565000 ;
        RECT 11.205000  0.085000 11.455000 0.565000 ;
        RECT 12.065000  0.085000 12.315000 0.565000 ;
        RECT 12.925000  0.085000 13.185000 0.565000 ;
        RECT 13.785000  0.085000 14.085000 0.565000 ;
      LAYER mcon ;
        RECT  0.145000 -0.085000  0.315000 0.085000 ;
        RECT  0.605000 -0.085000  0.775000 0.085000 ;
        RECT  1.065000 -0.085000  1.235000 0.085000 ;
        RECT  1.525000 -0.085000  1.695000 0.085000 ;
        RECT  1.985000 -0.085000  2.155000 0.085000 ;
        RECT  2.445000 -0.085000  2.615000 0.085000 ;
        RECT  2.905000 -0.085000  3.075000 0.085000 ;
        RECT  3.365000 -0.085000  3.535000 0.085000 ;
        RECT  3.825000 -0.085000  3.995000 0.085000 ;
        RECT  4.285000 -0.085000  4.455000 0.085000 ;
        RECT  4.745000 -0.085000  4.915000 0.085000 ;
        RECT  5.205000 -0.085000  5.375000 0.085000 ;
        RECT  5.665000 -0.085000  5.835000 0.085000 ;
        RECT  6.125000 -0.085000  6.295000 0.085000 ;
        RECT  6.585000 -0.085000  6.755000 0.085000 ;
        RECT  7.045000 -0.085000  7.215000 0.085000 ;
        RECT  7.505000 -0.085000  7.675000 0.085000 ;
        RECT  7.965000 -0.085000  8.135000 0.085000 ;
        RECT  8.425000 -0.085000  8.595000 0.085000 ;
        RECT  8.885000 -0.085000  9.055000 0.085000 ;
        RECT  9.345000 -0.085000  9.515000 0.085000 ;
        RECT  9.805000 -0.085000  9.975000 0.085000 ;
        RECT 10.265000 -0.085000 10.435000 0.085000 ;
        RECT 10.725000 -0.085000 10.895000 0.085000 ;
        RECT 11.185000 -0.085000 11.355000 0.085000 ;
        RECT 11.645000 -0.085000 11.815000 0.085000 ;
        RECT 12.105000 -0.085000 12.275000 0.085000 ;
        RECT 12.565000 -0.085000 12.735000 0.085000 ;
        RECT 13.025000 -0.085000 13.195000 0.085000 ;
        RECT 13.485000 -0.085000 13.655000 0.085000 ;
        RECT 13.945000 -0.085000 14.115000 0.085000 ;
      LAYER met1 ;
        RECT 0.000000 -0.240000 14.260000 0.240000 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INOUT ;
    SHAPE ABUTMENT ;
    USE POWER ;
    PORT
      LAYER li1 ;
        RECT 0.000000 2.635000 14.260000 2.805000 ;
        RECT 0.130000 1.495000  0.535000 2.635000 ;
        RECT 3.435000 1.835000  3.685000 2.635000 ;
        RECT 4.195000 1.835000  4.525000 2.635000 ;
      LAYER mcon ;
        RECT  0.145000 2.635000  0.315000 2.805000 ;
        RECT  0.605000 2.635000  0.775000 2.805000 ;
        RECT  1.065000 2.635000  1.235000 2.805000 ;
        RECT  1.525000 2.635000  1.695000 2.805000 ;
        RECT  1.985000 2.635000  2.155000 2.805000 ;
        RECT  2.445000 2.635000  2.615000 2.805000 ;
        RECT  2.905000 2.635000  3.075000 2.805000 ;
        RECT  3.365000 2.635000  3.535000 2.805000 ;
        RECT  3.825000 2.635000  3.995000 2.805000 ;
        RECT  4.285000 2.635000  4.455000 2.805000 ;
        RECT  4.745000 2.635000  4.915000 2.805000 ;
        RECT  5.205000 2.635000  5.375000 2.805000 ;
        RECT  5.665000 2.635000  5.835000 2.805000 ;
        RECT  6.125000 2.635000  6.295000 2.805000 ;
        RECT  6.585000 2.635000  6.755000 2.805000 ;
        RECT  7.045000 2.635000  7.215000 2.805000 ;
        RECT  7.505000 2.635000  7.675000 2.805000 ;
        RECT  7.965000 2.635000  8.135000 2.805000 ;
        RECT  8.425000 2.635000  8.595000 2.805000 ;
        RECT  8.885000 2.635000  9.055000 2.805000 ;
        RECT  9.345000 2.635000  9.515000 2.805000 ;
        RECT  9.805000 2.635000  9.975000 2.805000 ;
        RECT 10.265000 2.635000 10.435000 2.805000 ;
        RECT 10.725000 2.635000 10.895000 2.805000 ;
        RECT 11.185000 2.635000 11.355000 2.805000 ;
        RECT 11.645000 2.635000 11.815000 2.805000 ;
        RECT 12.105000 2.635000 12.275000 2.805000 ;
        RECT 12.565000 2.635000 12.735000 2.805000 ;
        RECT 13.025000 2.635000 13.195000 2.805000 ;
        RECT 13.485000 2.635000 13.655000 2.805000 ;
        RECT 13.945000 2.635000 14.115000 2.805000 ;
      LAYER met1 ;
        RECT 0.000000 2.480000 14.260000 2.960000 ;
    END
  END VPWR
  OBS
    LAYER li1 ;
      RECT 0.705000 0.255000  1.035000 0.815000 ;
      RECT 0.705000 1.575000  1.035000 2.465000 ;
      RECT 0.785000 0.815000  1.035000 1.075000 ;
      RECT 0.785000 1.075000  2.265000 1.275000 ;
      RECT 0.785000 1.275000  1.035000 1.575000 ;
      RECT 1.205000 1.575000  1.585000 2.295000 ;
      RECT 1.205000 2.295000  3.265000 2.465000 ;
      RECT 1.675000 0.255000  2.005000 0.725000 ;
      RECT 1.675000 0.725000  4.525000 0.905000 ;
      RECT 1.755000 1.445000  2.765000 1.745000 ;
      RECT 1.755000 1.745000  1.925000 2.125000 ;
      RECT 2.095000 1.935000  2.425000 2.295000 ;
      RECT 2.435000 0.905000  3.095000 0.965000 ;
      RECT 2.435000 0.965000  2.765000 1.445000 ;
      RECT 2.515000 0.255000  2.845000 0.725000 ;
      RECT 2.595000 1.745000  2.765000 2.125000 ;
      RECT 2.935000 1.455000  4.975000 1.665000 ;
      RECT 2.935000 1.665000  3.265000 2.295000 ;
      RECT 3.355000 0.255000  3.685000 0.725000 ;
      RECT 3.855000 1.665000  4.025000 2.465000 ;
      RECT 4.195000 0.255000  4.525000 0.725000 ;
      RECT 4.695000 1.665000  4.975000 2.465000 ;
      RECT 5.145000 0.735000  5.460000 1.325000 ;
      RECT 5.655000 0.265000  5.880000 1.075000 ;
      RECT 5.655000 1.075000 12.750000 1.325000 ;
      RECT 5.655000 1.325000  5.845000 2.465000 ;
      RECT 6.490000 0.265000  6.740000 1.075000 ;
      RECT 6.515000 1.325000  6.705000 2.460000 ;
    LAYER mcon ;
      RECT 2.525000 0.765000 2.695000 0.935000 ;
      RECT 2.885000 0.765000 3.055000 0.935000 ;
      RECT 5.210000 0.765000 5.380000 0.935000 ;
    LAYER met1 ;
      RECT 2.465000 0.735000 3.115000 0.780000 ;
      RECT 2.465000 0.780000 5.440000 0.920000 ;
      RECT 2.465000 0.920000 3.115000 0.965000 ;
      RECT 5.150000 0.735000 5.440000 0.780000 ;
      RECT 5.150000 0.920000 5.440000 0.965000 ;
  END
END sky130_fd_sc_hd__lpflow_isobufsrckapwr_16
END LIBRARY
